// Generator : SpinalHDL v1.7.0    git head : eca519e78d4e6022e34911ec300a432ed9db8220
// Component : AES_ENGINE

`timescale 1ns/1ps 
module AES_ENGINE (
  input               io_engine_cmd_valid,
  output              io_engine_cmd_ready,
  input      [127:0]  io_engine_cmd_payload_key,
  input      [127:0]  io_engine_cmd_payload_block,
  input               io_engine_cmd_payload_enc,
  output              io_engine_rsp_valid,
  output     [127:0]  io_engine_rsp_payload_block,
  input               clk,
  input               reset
);

  reg        [127:0]  rndFuc_io_roundData;
  reg                 rndFuc_io_needMix;
  wire       [7:0]    _zz_CtrlState_keyRcon_port0;
  wire       [127:0]  rndFuc_io_result;
  reg                 CtrlState_enginRdy;
  reg                 CtrlState_ongoing;
  reg        [127:0]  CtrlState_nextrndKey;
  reg        [3:0]    CtrlState_rndCnt;
  reg        [127:0]  CtrlState_dataBuf;
  wire                CtrlState_lastRound;
  reg        [127:0]  CtrlState_currndKey;
  wire                io_engine_cmd_fire;
  wire                io_engine_cmd_fire_1;
  wire       [127:0]  _zz_CtrlState_nextrndKey;
  wire       [31:0]   _zz_CtrlState_nextrndKey_1;
  wire       [31:0]   _zz_CtrlState_nextrndKey_2;
  wire       [31:0]   _zz_CtrlState_nextrndKey_3;
  wire       [31:0]   _zz_CtrlState_nextrndKey_4;
  wire       [31:0]   _zz_CtrlState_nextrndKey_5;
  reg        [31:0]   _zz_CtrlState_nextrndKey_6;
  wire       [7:0]    _zz_CtrlState_nextrndKey_7;
  reg        [7:0]    _zz_CtrlState_nextrndKey_8;
  wire       [7:0]    _zz_CtrlState_nextrndKey_9;
  reg        [7:0]    _zz_CtrlState_nextrndKey_10;
  wire       [7:0]    _zz_CtrlState_nextrndKey_11;
  reg        [7:0]    _zz_CtrlState_nextrndKey_12;
  wire       [3:0]    _zz_CtrlState_nextrndKey_13;
  wire       [3:0]    _zz_CtrlState_nextrndKey_14;
  wire       [3:0]    _zz_CtrlState_nextrndKey_15;
  reg        [3:0]    _zz_CtrlState_nextrndKey_16;
  reg        [3:0]    _zz_CtrlState_nextrndKey_17;
  wire       [1:0]    _zz_CtrlState_nextrndKey_18;
  wire       [1:0]    _zz_CtrlState_nextrndKey_19;
  wire       [1:0]    _zz_CtrlState_nextrndKey_20;
  wire       [1:0]    _zz_CtrlState_nextrndKey_21;
  wire       [1:0]    _zz_CtrlState_nextrndKey_22;
  wire       [1:0]    _zz_CtrlState_nextrndKey_23;
  wire       [1:0]    _zz_CtrlState_nextrndKey_24;
  wire                _zz_CtrlState_nextrndKey_25;
  reg        [1:0]    _zz_CtrlState_nextrndKey_26;
  wire       [1:0]    _zz_CtrlState_nextrndKey_27;
  reg        [1:0]    _zz_CtrlState_nextrndKey_28;
  wire                _zz_CtrlState_nextrndKey_29;
  reg        [1:0]    _zz_CtrlState_nextrndKey_30;
  wire                _zz_CtrlState_nextrndKey_31;
  reg        [1:0]    _zz_CtrlState_nextrndKey_32;
  wire       [3:0]    _zz_CtrlState_nextrndKey_33;
  wire       [3:0]    _zz_CtrlState_nextrndKey_34;
  reg        [3:0]    _zz_CtrlState_nextrndKey_35;
  wire       [1:0]    _zz_CtrlState_nextrndKey_36;
  wire       [1:0]    _zz_CtrlState_nextrndKey_37;
  wire       [1:0]    _zz_CtrlState_nextrndKey_38;
  reg        [1:0]    _zz_CtrlState_nextrndKey_39;
  wire                _zz_CtrlState_nextrndKey_40;
  reg        [1:0]    _zz_CtrlState_nextrndKey_41;
  wire       [1:0]    _zz_CtrlState_nextrndKey_42;
  wire       [1:0]    _zz_CtrlState_nextrndKey_43;
  reg        [1:0]    _zz_CtrlState_nextrndKey_44;
  wire                _zz_CtrlState_nextrndKey_45;
  reg        [1:0]    _zz_CtrlState_nextrndKey_46;
  wire                _zz_CtrlState_nextrndKey_47;
  reg        [1:0]    _zz_CtrlState_nextrndKey_48;
  reg        [3:0]    _zz_CtrlState_nextrndKey_49;
  wire       [1:0]    _zz_CtrlState_nextrndKey_50;
  wire       [1:0]    _zz_CtrlState_nextrndKey_51;
  wire       [1:0]    _zz_CtrlState_nextrndKey_52;
  wire       [1:0]    _zz_CtrlState_nextrndKey_53;
  wire       [1:0]    _zz_CtrlState_nextrndKey_54;
  wire       [1:0]    _zz_CtrlState_nextrndKey_55;
  wire       [1:0]    _zz_CtrlState_nextrndKey_56;
  wire                _zz_CtrlState_nextrndKey_57;
  reg        [1:0]    _zz_CtrlState_nextrndKey_58;
  wire       [1:0]    _zz_CtrlState_nextrndKey_59;
  reg        [1:0]    _zz_CtrlState_nextrndKey_60;
  wire                _zz_CtrlState_nextrndKey_61;
  reg        [1:0]    _zz_CtrlState_nextrndKey_62;
  wire                _zz_CtrlState_nextrndKey_63;
  reg        [1:0]    _zz_CtrlState_nextrndKey_64;
  reg        [3:0]    _zz_CtrlState_nextrndKey_65;
  wire       [1:0]    _zz_CtrlState_nextrndKey_66;
  wire       [1:0]    _zz_CtrlState_nextrndKey_67;
  wire       [1:0]    _zz_CtrlState_nextrndKey_68;
  wire       [1:0]    _zz_CtrlState_nextrndKey_69;
  wire       [1:0]    _zz_CtrlState_nextrndKey_70;
  wire       [1:0]    _zz_CtrlState_nextrndKey_71;
  wire       [1:0]    _zz_CtrlState_nextrndKey_72;
  wire                _zz_CtrlState_nextrndKey_73;
  reg        [1:0]    _zz_CtrlState_nextrndKey_74;
  wire       [1:0]    _zz_CtrlState_nextrndKey_75;
  reg        [1:0]    _zz_CtrlState_nextrndKey_76;
  wire                _zz_CtrlState_nextrndKey_77;
  reg        [1:0]    _zz_CtrlState_nextrndKey_78;
  wire                _zz_CtrlState_nextrndKey_79;
  reg        [1:0]    _zz_CtrlState_nextrndKey_80;
  wire       [7:0]    _zz_CtrlState_nextrndKey_81;
  reg        [7:0]    _zz_CtrlState_nextrndKey_82;
  wire       [7:0]    _zz_CtrlState_nextrndKey_83;
  reg        [7:0]    _zz_CtrlState_nextrndKey_84;
  wire       [7:0]    _zz_CtrlState_nextrndKey_85;
  reg        [7:0]    _zz_CtrlState_nextrndKey_86;
  wire       [7:0]    _zz_CtrlState_nextrndKey_87;
  reg        [7:0]    _zz_CtrlState_nextrndKey_88;
  wire       [3:0]    _zz_CtrlState_nextrndKey_89;
  wire       [3:0]    _zz_CtrlState_nextrndKey_90;
  wire       [3:0]    _zz_CtrlState_nextrndKey_91;
  reg        [3:0]    _zz_CtrlState_nextrndKey_92;
  reg        [3:0]    _zz_CtrlState_nextrndKey_93;
  wire       [1:0]    _zz_CtrlState_nextrndKey_94;
  wire       [1:0]    _zz_CtrlState_nextrndKey_95;
  wire       [1:0]    _zz_CtrlState_nextrndKey_96;
  wire       [1:0]    _zz_CtrlState_nextrndKey_97;
  wire       [1:0]    _zz_CtrlState_nextrndKey_98;
  wire       [1:0]    _zz_CtrlState_nextrndKey_99;
  wire       [1:0]    _zz_CtrlState_nextrndKey_100;
  wire                _zz_CtrlState_nextrndKey_101;
  reg        [1:0]    _zz_CtrlState_nextrndKey_102;
  wire       [1:0]    _zz_CtrlState_nextrndKey_103;
  reg        [1:0]    _zz_CtrlState_nextrndKey_104;
  wire                _zz_CtrlState_nextrndKey_105;
  reg        [1:0]    _zz_CtrlState_nextrndKey_106;
  wire                _zz_CtrlState_nextrndKey_107;
  reg        [1:0]    _zz_CtrlState_nextrndKey_108;
  wire       [3:0]    _zz_CtrlState_nextrndKey_109;
  wire       [3:0]    _zz_CtrlState_nextrndKey_110;
  reg        [3:0]    _zz_CtrlState_nextrndKey_111;
  wire       [1:0]    _zz_CtrlState_nextrndKey_112;
  wire       [1:0]    _zz_CtrlState_nextrndKey_113;
  wire       [1:0]    _zz_CtrlState_nextrndKey_114;
  reg        [1:0]    _zz_CtrlState_nextrndKey_115;
  wire                _zz_CtrlState_nextrndKey_116;
  reg        [1:0]    _zz_CtrlState_nextrndKey_117;
  wire       [1:0]    _zz_CtrlState_nextrndKey_118;
  wire       [1:0]    _zz_CtrlState_nextrndKey_119;
  reg        [1:0]    _zz_CtrlState_nextrndKey_120;
  wire                _zz_CtrlState_nextrndKey_121;
  reg        [1:0]    _zz_CtrlState_nextrndKey_122;
  wire                _zz_CtrlState_nextrndKey_123;
  reg        [1:0]    _zz_CtrlState_nextrndKey_124;
  reg        [3:0]    _zz_CtrlState_nextrndKey_125;
  wire       [1:0]    _zz_CtrlState_nextrndKey_126;
  wire       [1:0]    _zz_CtrlState_nextrndKey_127;
  wire       [1:0]    _zz_CtrlState_nextrndKey_128;
  wire       [1:0]    _zz_CtrlState_nextrndKey_129;
  wire       [1:0]    _zz_CtrlState_nextrndKey_130;
  wire       [1:0]    _zz_CtrlState_nextrndKey_131;
  wire       [1:0]    _zz_CtrlState_nextrndKey_132;
  wire                _zz_CtrlState_nextrndKey_133;
  reg        [1:0]    _zz_CtrlState_nextrndKey_134;
  wire       [1:0]    _zz_CtrlState_nextrndKey_135;
  reg        [1:0]    _zz_CtrlState_nextrndKey_136;
  wire                _zz_CtrlState_nextrndKey_137;
  reg        [1:0]    _zz_CtrlState_nextrndKey_138;
  wire                _zz_CtrlState_nextrndKey_139;
  reg        [1:0]    _zz_CtrlState_nextrndKey_140;
  reg        [3:0]    _zz_CtrlState_nextrndKey_141;
  wire       [1:0]    _zz_CtrlState_nextrndKey_142;
  wire       [1:0]    _zz_CtrlState_nextrndKey_143;
  wire       [1:0]    _zz_CtrlState_nextrndKey_144;
  wire       [1:0]    _zz_CtrlState_nextrndKey_145;
  wire       [1:0]    _zz_CtrlState_nextrndKey_146;
  wire       [1:0]    _zz_CtrlState_nextrndKey_147;
  wire       [1:0]    _zz_CtrlState_nextrndKey_148;
  wire                _zz_CtrlState_nextrndKey_149;
  reg        [1:0]    _zz_CtrlState_nextrndKey_150;
  wire       [1:0]    _zz_CtrlState_nextrndKey_151;
  reg        [1:0]    _zz_CtrlState_nextrndKey_152;
  wire                _zz_CtrlState_nextrndKey_153;
  reg        [1:0]    _zz_CtrlState_nextrndKey_154;
  wire                _zz_CtrlState_nextrndKey_155;
  reg        [1:0]    _zz_CtrlState_nextrndKey_156;
  wire       [7:0]    _zz_CtrlState_nextrndKey_157;
  reg        [7:0]    _zz_CtrlState_nextrndKey_158;
  wire       [7:0]    _zz_CtrlState_nextrndKey_159;
  reg        [7:0]    _zz_CtrlState_nextrndKey_160;
  wire       [7:0]    _zz_CtrlState_nextrndKey_161;
  reg        [7:0]    _zz_CtrlState_nextrndKey_162;
  wire       [7:0]    _zz_CtrlState_nextrndKey_163;
  reg        [7:0]    _zz_CtrlState_nextrndKey_164;
  wire       [3:0]    _zz_CtrlState_nextrndKey_165;
  wire       [3:0]    _zz_CtrlState_nextrndKey_166;
  wire       [3:0]    _zz_CtrlState_nextrndKey_167;
  reg        [3:0]    _zz_CtrlState_nextrndKey_168;
  reg        [3:0]    _zz_CtrlState_nextrndKey_169;
  wire       [1:0]    _zz_CtrlState_nextrndKey_170;
  wire       [1:0]    _zz_CtrlState_nextrndKey_171;
  wire       [1:0]    _zz_CtrlState_nextrndKey_172;
  wire       [1:0]    _zz_CtrlState_nextrndKey_173;
  wire       [1:0]    _zz_CtrlState_nextrndKey_174;
  wire       [1:0]    _zz_CtrlState_nextrndKey_175;
  wire       [1:0]    _zz_CtrlState_nextrndKey_176;
  wire                _zz_CtrlState_nextrndKey_177;
  reg        [1:0]    _zz_CtrlState_nextrndKey_178;
  wire       [1:0]    _zz_CtrlState_nextrndKey_179;
  reg        [1:0]    _zz_CtrlState_nextrndKey_180;
  wire                _zz_CtrlState_nextrndKey_181;
  reg        [1:0]    _zz_CtrlState_nextrndKey_182;
  wire                _zz_CtrlState_nextrndKey_183;
  reg        [1:0]    _zz_CtrlState_nextrndKey_184;
  wire       [3:0]    _zz_CtrlState_nextrndKey_185;
  wire       [3:0]    _zz_CtrlState_nextrndKey_186;
  reg        [3:0]    _zz_CtrlState_nextrndKey_187;
  wire       [1:0]    _zz_CtrlState_nextrndKey_188;
  wire       [1:0]    _zz_CtrlState_nextrndKey_189;
  wire       [1:0]    _zz_CtrlState_nextrndKey_190;
  reg        [1:0]    _zz_CtrlState_nextrndKey_191;
  wire                _zz_CtrlState_nextrndKey_192;
  reg        [1:0]    _zz_CtrlState_nextrndKey_193;
  wire       [1:0]    _zz_CtrlState_nextrndKey_194;
  wire       [1:0]    _zz_CtrlState_nextrndKey_195;
  reg        [1:0]    _zz_CtrlState_nextrndKey_196;
  wire                _zz_CtrlState_nextrndKey_197;
  reg        [1:0]    _zz_CtrlState_nextrndKey_198;
  wire                _zz_CtrlState_nextrndKey_199;
  reg        [1:0]    _zz_CtrlState_nextrndKey_200;
  reg        [3:0]    _zz_CtrlState_nextrndKey_201;
  wire       [1:0]    _zz_CtrlState_nextrndKey_202;
  wire       [1:0]    _zz_CtrlState_nextrndKey_203;
  wire       [1:0]    _zz_CtrlState_nextrndKey_204;
  wire       [1:0]    _zz_CtrlState_nextrndKey_205;
  wire       [1:0]    _zz_CtrlState_nextrndKey_206;
  wire       [1:0]    _zz_CtrlState_nextrndKey_207;
  wire       [1:0]    _zz_CtrlState_nextrndKey_208;
  wire                _zz_CtrlState_nextrndKey_209;
  reg        [1:0]    _zz_CtrlState_nextrndKey_210;
  wire       [1:0]    _zz_CtrlState_nextrndKey_211;
  reg        [1:0]    _zz_CtrlState_nextrndKey_212;
  wire                _zz_CtrlState_nextrndKey_213;
  reg        [1:0]    _zz_CtrlState_nextrndKey_214;
  wire                _zz_CtrlState_nextrndKey_215;
  reg        [1:0]    _zz_CtrlState_nextrndKey_216;
  reg        [3:0]    _zz_CtrlState_nextrndKey_217;
  wire       [1:0]    _zz_CtrlState_nextrndKey_218;
  wire       [1:0]    _zz_CtrlState_nextrndKey_219;
  wire       [1:0]    _zz_CtrlState_nextrndKey_220;
  wire       [1:0]    _zz_CtrlState_nextrndKey_221;
  wire       [1:0]    _zz_CtrlState_nextrndKey_222;
  wire       [1:0]    _zz_CtrlState_nextrndKey_223;
  wire       [1:0]    _zz_CtrlState_nextrndKey_224;
  wire                _zz_CtrlState_nextrndKey_225;
  reg        [1:0]    _zz_CtrlState_nextrndKey_226;
  wire       [1:0]    _zz_CtrlState_nextrndKey_227;
  reg        [1:0]    _zz_CtrlState_nextrndKey_228;
  wire                _zz_CtrlState_nextrndKey_229;
  reg        [1:0]    _zz_CtrlState_nextrndKey_230;
  wire                _zz_CtrlState_nextrndKey_231;
  reg        [1:0]    _zz_CtrlState_nextrndKey_232;
  wire       [7:0]    _zz_CtrlState_nextrndKey_233;
  reg        [7:0]    _zz_CtrlState_nextrndKey_234;
  wire       [7:0]    _zz_CtrlState_nextrndKey_235;
  reg        [7:0]    _zz_CtrlState_nextrndKey_236;
  wire       [7:0]    _zz_CtrlState_nextrndKey_237;
  reg        [7:0]    _zz_CtrlState_nextrndKey_238;
  wire       [7:0]    _zz_CtrlState_nextrndKey_239;
  reg        [7:0]    _zz_CtrlState_nextrndKey_240;
  wire       [3:0]    _zz_CtrlState_nextrndKey_241;
  wire       [3:0]    _zz_CtrlState_nextrndKey_242;
  wire       [3:0]    _zz_CtrlState_nextrndKey_243;
  reg        [3:0]    _zz_CtrlState_nextrndKey_244;
  reg        [3:0]    _zz_CtrlState_nextrndKey_245;
  wire       [1:0]    _zz_CtrlState_nextrndKey_246;
  wire       [1:0]    _zz_CtrlState_nextrndKey_247;
  wire       [1:0]    _zz_CtrlState_nextrndKey_248;
  wire       [1:0]    _zz_CtrlState_nextrndKey_249;
  wire       [1:0]    _zz_CtrlState_nextrndKey_250;
  wire       [1:0]    _zz_CtrlState_nextrndKey_251;
  wire       [1:0]    _zz_CtrlState_nextrndKey_252;
  wire                _zz_CtrlState_nextrndKey_253;
  reg        [1:0]    _zz_CtrlState_nextrndKey_254;
  wire       [1:0]    _zz_CtrlState_nextrndKey_255;
  reg        [1:0]    _zz_CtrlState_nextrndKey_256;
  wire                _zz_CtrlState_nextrndKey_257;
  reg        [1:0]    _zz_CtrlState_nextrndKey_258;
  wire                _zz_CtrlState_nextrndKey_259;
  reg        [1:0]    _zz_CtrlState_nextrndKey_260;
  wire       [3:0]    _zz_CtrlState_nextrndKey_261;
  wire       [3:0]    _zz_CtrlState_nextrndKey_262;
  reg        [3:0]    _zz_CtrlState_nextrndKey_263;
  wire       [1:0]    _zz_CtrlState_nextrndKey_264;
  wire       [1:0]    _zz_CtrlState_nextrndKey_265;
  wire       [1:0]    _zz_CtrlState_nextrndKey_266;
  reg        [1:0]    _zz_CtrlState_nextrndKey_267;
  wire                _zz_CtrlState_nextrndKey_268;
  reg        [1:0]    _zz_CtrlState_nextrndKey_269;
  wire       [1:0]    _zz_CtrlState_nextrndKey_270;
  wire       [1:0]    _zz_CtrlState_nextrndKey_271;
  reg        [1:0]    _zz_CtrlState_nextrndKey_272;
  wire                _zz_CtrlState_nextrndKey_273;
  reg        [1:0]    _zz_CtrlState_nextrndKey_274;
  wire                _zz_CtrlState_nextrndKey_275;
  reg        [1:0]    _zz_CtrlState_nextrndKey_276;
  reg        [3:0]    _zz_CtrlState_nextrndKey_277;
  wire       [1:0]    _zz_CtrlState_nextrndKey_278;
  wire       [1:0]    _zz_CtrlState_nextrndKey_279;
  wire       [1:0]    _zz_CtrlState_nextrndKey_280;
  wire       [1:0]    _zz_CtrlState_nextrndKey_281;
  wire       [1:0]    _zz_CtrlState_nextrndKey_282;
  wire       [1:0]    _zz_CtrlState_nextrndKey_283;
  wire       [1:0]    _zz_CtrlState_nextrndKey_284;
  wire                _zz_CtrlState_nextrndKey_285;
  reg        [1:0]    _zz_CtrlState_nextrndKey_286;
  wire       [1:0]    _zz_CtrlState_nextrndKey_287;
  reg        [1:0]    _zz_CtrlState_nextrndKey_288;
  wire                _zz_CtrlState_nextrndKey_289;
  reg        [1:0]    _zz_CtrlState_nextrndKey_290;
  wire                _zz_CtrlState_nextrndKey_291;
  reg        [1:0]    _zz_CtrlState_nextrndKey_292;
  reg        [3:0]    _zz_CtrlState_nextrndKey_293;
  wire       [1:0]    _zz_CtrlState_nextrndKey_294;
  wire       [1:0]    _zz_CtrlState_nextrndKey_295;
  wire       [1:0]    _zz_CtrlState_nextrndKey_296;
  wire       [1:0]    _zz_CtrlState_nextrndKey_297;
  wire       [1:0]    _zz_CtrlState_nextrndKey_298;
  wire       [1:0]    _zz_CtrlState_nextrndKey_299;
  wire       [1:0]    _zz_CtrlState_nextrndKey_300;
  wire                _zz_CtrlState_nextrndKey_301;
  reg        [1:0]    _zz_CtrlState_nextrndKey_302;
  wire       [1:0]    _zz_CtrlState_nextrndKey_303;
  reg        [1:0]    _zz_CtrlState_nextrndKey_304;
  wire                _zz_CtrlState_nextrndKey_305;
  reg        [1:0]    _zz_CtrlState_nextrndKey_306;
  wire                _zz_CtrlState_nextrndKey_307;
  reg        [1:0]    _zz_CtrlState_nextrndKey_308;
  wire       [7:0]    _zz_CtrlState_nextrndKey_309;
  reg        [7:0]    _zz_CtrlState_nextrndKey_310;
  wire       [127:0]  _zz_CtrlState_nextrndKey_311;
  wire       [3:0]    _zz_CtrlState_nextrndKey_312;
  wire       [31:0]   _zz_CtrlState_nextrndKey_313;
  wire       [31:0]   _zz_CtrlState_nextrndKey_314;
  wire       [31:0]   _zz_CtrlState_nextrndKey_315;
  wire       [31:0]   _zz_CtrlState_nextrndKey_316;
  wire       [31:0]   _zz_CtrlState_nextrndKey_317;
  reg        [31:0]   _zz_CtrlState_nextrndKey_318;
  wire       [7:0]    _zz_CtrlState_nextrndKey_319;
  reg        [7:0]    _zz_CtrlState_nextrndKey_320;
  wire       [7:0]    _zz_CtrlState_nextrndKey_321;
  reg        [7:0]    _zz_CtrlState_nextrndKey_322;
  wire       [7:0]    _zz_CtrlState_nextrndKey_323;
  reg        [7:0]    _zz_CtrlState_nextrndKey_324;
  wire       [3:0]    _zz_CtrlState_nextrndKey_325;
  wire       [3:0]    _zz_CtrlState_nextrndKey_326;
  wire       [3:0]    _zz_CtrlState_nextrndKey_327;
  reg        [3:0]    _zz_CtrlState_nextrndKey_328;
  reg        [3:0]    _zz_CtrlState_nextrndKey_329;
  wire       [1:0]    _zz_CtrlState_nextrndKey_330;
  wire       [1:0]    _zz_CtrlState_nextrndKey_331;
  wire       [1:0]    _zz_CtrlState_nextrndKey_332;
  wire       [1:0]    _zz_CtrlState_nextrndKey_333;
  wire       [1:0]    _zz_CtrlState_nextrndKey_334;
  wire       [1:0]    _zz_CtrlState_nextrndKey_335;
  wire       [1:0]    _zz_CtrlState_nextrndKey_336;
  wire                _zz_CtrlState_nextrndKey_337;
  reg        [1:0]    _zz_CtrlState_nextrndKey_338;
  wire       [1:0]    _zz_CtrlState_nextrndKey_339;
  reg        [1:0]    _zz_CtrlState_nextrndKey_340;
  wire                _zz_CtrlState_nextrndKey_341;
  reg        [1:0]    _zz_CtrlState_nextrndKey_342;
  wire                _zz_CtrlState_nextrndKey_343;
  reg        [1:0]    _zz_CtrlState_nextrndKey_344;
  wire       [3:0]    _zz_CtrlState_nextrndKey_345;
  wire       [3:0]    _zz_CtrlState_nextrndKey_346;
  reg        [3:0]    _zz_CtrlState_nextrndKey_347;
  wire       [1:0]    _zz_CtrlState_nextrndKey_348;
  wire       [1:0]    _zz_CtrlState_nextrndKey_349;
  wire       [1:0]    _zz_CtrlState_nextrndKey_350;
  reg        [1:0]    _zz_CtrlState_nextrndKey_351;
  wire                _zz_CtrlState_nextrndKey_352;
  reg        [1:0]    _zz_CtrlState_nextrndKey_353;
  wire       [1:0]    _zz_CtrlState_nextrndKey_354;
  wire       [1:0]    _zz_CtrlState_nextrndKey_355;
  reg        [1:0]    _zz_CtrlState_nextrndKey_356;
  wire                _zz_CtrlState_nextrndKey_357;
  reg        [1:0]    _zz_CtrlState_nextrndKey_358;
  wire                _zz_CtrlState_nextrndKey_359;
  reg        [1:0]    _zz_CtrlState_nextrndKey_360;
  reg        [3:0]    _zz_CtrlState_nextrndKey_361;
  wire       [1:0]    _zz_CtrlState_nextrndKey_362;
  wire       [1:0]    _zz_CtrlState_nextrndKey_363;
  wire       [1:0]    _zz_CtrlState_nextrndKey_364;
  wire       [1:0]    _zz_CtrlState_nextrndKey_365;
  wire       [1:0]    _zz_CtrlState_nextrndKey_366;
  wire       [1:0]    _zz_CtrlState_nextrndKey_367;
  wire       [1:0]    _zz_CtrlState_nextrndKey_368;
  wire                _zz_CtrlState_nextrndKey_369;
  reg        [1:0]    _zz_CtrlState_nextrndKey_370;
  wire       [1:0]    _zz_CtrlState_nextrndKey_371;
  reg        [1:0]    _zz_CtrlState_nextrndKey_372;
  wire                _zz_CtrlState_nextrndKey_373;
  reg        [1:0]    _zz_CtrlState_nextrndKey_374;
  wire                _zz_CtrlState_nextrndKey_375;
  reg        [1:0]    _zz_CtrlState_nextrndKey_376;
  reg        [3:0]    _zz_CtrlState_nextrndKey_377;
  wire       [1:0]    _zz_CtrlState_nextrndKey_378;
  wire       [1:0]    _zz_CtrlState_nextrndKey_379;
  wire       [1:0]    _zz_CtrlState_nextrndKey_380;
  wire       [1:0]    _zz_CtrlState_nextrndKey_381;
  wire       [1:0]    _zz_CtrlState_nextrndKey_382;
  wire       [1:0]    _zz_CtrlState_nextrndKey_383;
  wire       [1:0]    _zz_CtrlState_nextrndKey_384;
  wire                _zz_CtrlState_nextrndKey_385;
  reg        [1:0]    _zz_CtrlState_nextrndKey_386;
  wire       [1:0]    _zz_CtrlState_nextrndKey_387;
  reg        [1:0]    _zz_CtrlState_nextrndKey_388;
  wire                _zz_CtrlState_nextrndKey_389;
  reg        [1:0]    _zz_CtrlState_nextrndKey_390;
  wire                _zz_CtrlState_nextrndKey_391;
  reg        [1:0]    _zz_CtrlState_nextrndKey_392;
  wire       [7:0]    _zz_CtrlState_nextrndKey_393;
  reg        [7:0]    _zz_CtrlState_nextrndKey_394;
  wire       [7:0]    _zz_CtrlState_nextrndKey_395;
  reg        [7:0]    _zz_CtrlState_nextrndKey_396;
  wire       [7:0]    _zz_CtrlState_nextrndKey_397;
  reg        [7:0]    _zz_CtrlState_nextrndKey_398;
  wire       [7:0]    _zz_CtrlState_nextrndKey_399;
  reg        [7:0]    _zz_CtrlState_nextrndKey_400;
  wire       [3:0]    _zz_CtrlState_nextrndKey_401;
  wire       [3:0]    _zz_CtrlState_nextrndKey_402;
  wire       [3:0]    _zz_CtrlState_nextrndKey_403;
  reg        [3:0]    _zz_CtrlState_nextrndKey_404;
  reg        [3:0]    _zz_CtrlState_nextrndKey_405;
  wire       [1:0]    _zz_CtrlState_nextrndKey_406;
  wire       [1:0]    _zz_CtrlState_nextrndKey_407;
  wire       [1:0]    _zz_CtrlState_nextrndKey_408;
  wire       [1:0]    _zz_CtrlState_nextrndKey_409;
  wire       [1:0]    _zz_CtrlState_nextrndKey_410;
  wire       [1:0]    _zz_CtrlState_nextrndKey_411;
  wire       [1:0]    _zz_CtrlState_nextrndKey_412;
  wire                _zz_CtrlState_nextrndKey_413;
  reg        [1:0]    _zz_CtrlState_nextrndKey_414;
  wire       [1:0]    _zz_CtrlState_nextrndKey_415;
  reg        [1:0]    _zz_CtrlState_nextrndKey_416;
  wire                _zz_CtrlState_nextrndKey_417;
  reg        [1:0]    _zz_CtrlState_nextrndKey_418;
  wire                _zz_CtrlState_nextrndKey_419;
  reg        [1:0]    _zz_CtrlState_nextrndKey_420;
  wire       [3:0]    _zz_CtrlState_nextrndKey_421;
  wire       [3:0]    _zz_CtrlState_nextrndKey_422;
  reg        [3:0]    _zz_CtrlState_nextrndKey_423;
  wire       [1:0]    _zz_CtrlState_nextrndKey_424;
  wire       [1:0]    _zz_CtrlState_nextrndKey_425;
  wire       [1:0]    _zz_CtrlState_nextrndKey_426;
  reg        [1:0]    _zz_CtrlState_nextrndKey_427;
  wire                _zz_CtrlState_nextrndKey_428;
  reg        [1:0]    _zz_CtrlState_nextrndKey_429;
  wire       [1:0]    _zz_CtrlState_nextrndKey_430;
  wire       [1:0]    _zz_CtrlState_nextrndKey_431;
  reg        [1:0]    _zz_CtrlState_nextrndKey_432;
  wire                _zz_CtrlState_nextrndKey_433;
  reg        [1:0]    _zz_CtrlState_nextrndKey_434;
  wire                _zz_CtrlState_nextrndKey_435;
  reg        [1:0]    _zz_CtrlState_nextrndKey_436;
  reg        [3:0]    _zz_CtrlState_nextrndKey_437;
  wire       [1:0]    _zz_CtrlState_nextrndKey_438;
  wire       [1:0]    _zz_CtrlState_nextrndKey_439;
  wire       [1:0]    _zz_CtrlState_nextrndKey_440;
  wire       [1:0]    _zz_CtrlState_nextrndKey_441;
  wire       [1:0]    _zz_CtrlState_nextrndKey_442;
  wire       [1:0]    _zz_CtrlState_nextrndKey_443;
  wire       [1:0]    _zz_CtrlState_nextrndKey_444;
  wire                _zz_CtrlState_nextrndKey_445;
  reg        [1:0]    _zz_CtrlState_nextrndKey_446;
  wire       [1:0]    _zz_CtrlState_nextrndKey_447;
  reg        [1:0]    _zz_CtrlState_nextrndKey_448;
  wire                _zz_CtrlState_nextrndKey_449;
  reg        [1:0]    _zz_CtrlState_nextrndKey_450;
  wire                _zz_CtrlState_nextrndKey_451;
  reg        [1:0]    _zz_CtrlState_nextrndKey_452;
  reg        [3:0]    _zz_CtrlState_nextrndKey_453;
  wire       [1:0]    _zz_CtrlState_nextrndKey_454;
  wire       [1:0]    _zz_CtrlState_nextrndKey_455;
  wire       [1:0]    _zz_CtrlState_nextrndKey_456;
  wire       [1:0]    _zz_CtrlState_nextrndKey_457;
  wire       [1:0]    _zz_CtrlState_nextrndKey_458;
  wire       [1:0]    _zz_CtrlState_nextrndKey_459;
  wire       [1:0]    _zz_CtrlState_nextrndKey_460;
  wire                _zz_CtrlState_nextrndKey_461;
  reg        [1:0]    _zz_CtrlState_nextrndKey_462;
  wire       [1:0]    _zz_CtrlState_nextrndKey_463;
  reg        [1:0]    _zz_CtrlState_nextrndKey_464;
  wire                _zz_CtrlState_nextrndKey_465;
  reg        [1:0]    _zz_CtrlState_nextrndKey_466;
  wire                _zz_CtrlState_nextrndKey_467;
  reg        [1:0]    _zz_CtrlState_nextrndKey_468;
  wire       [7:0]    _zz_CtrlState_nextrndKey_469;
  reg        [7:0]    _zz_CtrlState_nextrndKey_470;
  wire       [7:0]    _zz_CtrlState_nextrndKey_471;
  reg        [7:0]    _zz_CtrlState_nextrndKey_472;
  wire       [7:0]    _zz_CtrlState_nextrndKey_473;
  reg        [7:0]    _zz_CtrlState_nextrndKey_474;
  wire       [7:0]    _zz_CtrlState_nextrndKey_475;
  reg        [7:0]    _zz_CtrlState_nextrndKey_476;
  wire       [3:0]    _zz_CtrlState_nextrndKey_477;
  wire       [3:0]    _zz_CtrlState_nextrndKey_478;
  wire       [3:0]    _zz_CtrlState_nextrndKey_479;
  reg        [3:0]    _zz_CtrlState_nextrndKey_480;
  reg        [3:0]    _zz_CtrlState_nextrndKey_481;
  wire       [1:0]    _zz_CtrlState_nextrndKey_482;
  wire       [1:0]    _zz_CtrlState_nextrndKey_483;
  wire       [1:0]    _zz_CtrlState_nextrndKey_484;
  wire       [1:0]    _zz_CtrlState_nextrndKey_485;
  wire       [1:0]    _zz_CtrlState_nextrndKey_486;
  wire       [1:0]    _zz_CtrlState_nextrndKey_487;
  wire       [1:0]    _zz_CtrlState_nextrndKey_488;
  wire                _zz_CtrlState_nextrndKey_489;
  reg        [1:0]    _zz_CtrlState_nextrndKey_490;
  wire       [1:0]    _zz_CtrlState_nextrndKey_491;
  reg        [1:0]    _zz_CtrlState_nextrndKey_492;
  wire                _zz_CtrlState_nextrndKey_493;
  reg        [1:0]    _zz_CtrlState_nextrndKey_494;
  wire                _zz_CtrlState_nextrndKey_495;
  reg        [1:0]    _zz_CtrlState_nextrndKey_496;
  wire       [3:0]    _zz_CtrlState_nextrndKey_497;
  wire       [3:0]    _zz_CtrlState_nextrndKey_498;
  reg        [3:0]    _zz_CtrlState_nextrndKey_499;
  wire       [1:0]    _zz_CtrlState_nextrndKey_500;
  wire       [1:0]    _zz_CtrlState_nextrndKey_501;
  wire       [1:0]    _zz_CtrlState_nextrndKey_502;
  reg        [1:0]    _zz_CtrlState_nextrndKey_503;
  wire                _zz_CtrlState_nextrndKey_504;
  reg        [1:0]    _zz_CtrlState_nextrndKey_505;
  wire       [1:0]    _zz_CtrlState_nextrndKey_506;
  wire       [1:0]    _zz_CtrlState_nextrndKey_507;
  reg        [1:0]    _zz_CtrlState_nextrndKey_508;
  wire                _zz_CtrlState_nextrndKey_509;
  reg        [1:0]    _zz_CtrlState_nextrndKey_510;
  wire                _zz_CtrlState_nextrndKey_511;
  reg        [1:0]    _zz_CtrlState_nextrndKey_512;
  reg        [3:0]    _zz_CtrlState_nextrndKey_513;
  wire       [1:0]    _zz_CtrlState_nextrndKey_514;
  wire       [1:0]    _zz_CtrlState_nextrndKey_515;
  wire       [1:0]    _zz_CtrlState_nextrndKey_516;
  wire       [1:0]    _zz_CtrlState_nextrndKey_517;
  wire       [1:0]    _zz_CtrlState_nextrndKey_518;
  wire       [1:0]    _zz_CtrlState_nextrndKey_519;
  wire       [1:0]    _zz_CtrlState_nextrndKey_520;
  wire                _zz_CtrlState_nextrndKey_521;
  reg        [1:0]    _zz_CtrlState_nextrndKey_522;
  wire       [1:0]    _zz_CtrlState_nextrndKey_523;
  reg        [1:0]    _zz_CtrlState_nextrndKey_524;
  wire                _zz_CtrlState_nextrndKey_525;
  reg        [1:0]    _zz_CtrlState_nextrndKey_526;
  wire                _zz_CtrlState_nextrndKey_527;
  reg        [1:0]    _zz_CtrlState_nextrndKey_528;
  reg        [3:0]    _zz_CtrlState_nextrndKey_529;
  wire       [1:0]    _zz_CtrlState_nextrndKey_530;
  wire       [1:0]    _zz_CtrlState_nextrndKey_531;
  wire       [1:0]    _zz_CtrlState_nextrndKey_532;
  wire       [1:0]    _zz_CtrlState_nextrndKey_533;
  wire       [1:0]    _zz_CtrlState_nextrndKey_534;
  wire       [1:0]    _zz_CtrlState_nextrndKey_535;
  wire       [1:0]    _zz_CtrlState_nextrndKey_536;
  wire                _zz_CtrlState_nextrndKey_537;
  reg        [1:0]    _zz_CtrlState_nextrndKey_538;
  wire       [1:0]    _zz_CtrlState_nextrndKey_539;
  reg        [1:0]    _zz_CtrlState_nextrndKey_540;
  wire                _zz_CtrlState_nextrndKey_541;
  reg        [1:0]    _zz_CtrlState_nextrndKey_542;
  wire                _zz_CtrlState_nextrndKey_543;
  reg        [1:0]    _zz_CtrlState_nextrndKey_544;
  wire       [7:0]    _zz_CtrlState_nextrndKey_545;
  reg        [7:0]    _zz_CtrlState_nextrndKey_546;
  wire       [7:0]    _zz_CtrlState_nextrndKey_547;
  reg        [7:0]    _zz_CtrlState_nextrndKey_548;
  wire       [7:0]    _zz_CtrlState_nextrndKey_549;
  reg        [7:0]    _zz_CtrlState_nextrndKey_550;
  wire       [7:0]    _zz_CtrlState_nextrndKey_551;
  reg        [7:0]    _zz_CtrlState_nextrndKey_552;
  wire       [3:0]    _zz_CtrlState_nextrndKey_553;
  wire       [3:0]    _zz_CtrlState_nextrndKey_554;
  wire       [3:0]    _zz_CtrlState_nextrndKey_555;
  reg        [3:0]    _zz_CtrlState_nextrndKey_556;
  reg        [3:0]    _zz_CtrlState_nextrndKey_557;
  wire       [1:0]    _zz_CtrlState_nextrndKey_558;
  wire       [1:0]    _zz_CtrlState_nextrndKey_559;
  wire       [1:0]    _zz_CtrlState_nextrndKey_560;
  wire       [1:0]    _zz_CtrlState_nextrndKey_561;
  wire       [1:0]    _zz_CtrlState_nextrndKey_562;
  wire       [1:0]    _zz_CtrlState_nextrndKey_563;
  wire       [1:0]    _zz_CtrlState_nextrndKey_564;
  wire                _zz_CtrlState_nextrndKey_565;
  reg        [1:0]    _zz_CtrlState_nextrndKey_566;
  wire       [1:0]    _zz_CtrlState_nextrndKey_567;
  reg        [1:0]    _zz_CtrlState_nextrndKey_568;
  wire                _zz_CtrlState_nextrndKey_569;
  reg        [1:0]    _zz_CtrlState_nextrndKey_570;
  wire                _zz_CtrlState_nextrndKey_571;
  reg        [1:0]    _zz_CtrlState_nextrndKey_572;
  wire       [3:0]    _zz_CtrlState_nextrndKey_573;
  wire       [3:0]    _zz_CtrlState_nextrndKey_574;
  reg        [3:0]    _zz_CtrlState_nextrndKey_575;
  wire       [1:0]    _zz_CtrlState_nextrndKey_576;
  wire       [1:0]    _zz_CtrlState_nextrndKey_577;
  wire       [1:0]    _zz_CtrlState_nextrndKey_578;
  reg        [1:0]    _zz_CtrlState_nextrndKey_579;
  wire                _zz_CtrlState_nextrndKey_580;
  reg        [1:0]    _zz_CtrlState_nextrndKey_581;
  wire       [1:0]    _zz_CtrlState_nextrndKey_582;
  wire       [1:0]    _zz_CtrlState_nextrndKey_583;
  reg        [1:0]    _zz_CtrlState_nextrndKey_584;
  wire                _zz_CtrlState_nextrndKey_585;
  reg        [1:0]    _zz_CtrlState_nextrndKey_586;
  wire                _zz_CtrlState_nextrndKey_587;
  reg        [1:0]    _zz_CtrlState_nextrndKey_588;
  reg        [3:0]    _zz_CtrlState_nextrndKey_589;
  wire       [1:0]    _zz_CtrlState_nextrndKey_590;
  wire       [1:0]    _zz_CtrlState_nextrndKey_591;
  wire       [1:0]    _zz_CtrlState_nextrndKey_592;
  wire       [1:0]    _zz_CtrlState_nextrndKey_593;
  wire       [1:0]    _zz_CtrlState_nextrndKey_594;
  wire       [1:0]    _zz_CtrlState_nextrndKey_595;
  wire       [1:0]    _zz_CtrlState_nextrndKey_596;
  wire                _zz_CtrlState_nextrndKey_597;
  reg        [1:0]    _zz_CtrlState_nextrndKey_598;
  wire       [1:0]    _zz_CtrlState_nextrndKey_599;
  reg        [1:0]    _zz_CtrlState_nextrndKey_600;
  wire                _zz_CtrlState_nextrndKey_601;
  reg        [1:0]    _zz_CtrlState_nextrndKey_602;
  wire                _zz_CtrlState_nextrndKey_603;
  reg        [1:0]    _zz_CtrlState_nextrndKey_604;
  reg        [3:0]    _zz_CtrlState_nextrndKey_605;
  wire       [1:0]    _zz_CtrlState_nextrndKey_606;
  wire       [1:0]    _zz_CtrlState_nextrndKey_607;
  wire       [1:0]    _zz_CtrlState_nextrndKey_608;
  wire       [1:0]    _zz_CtrlState_nextrndKey_609;
  wire       [1:0]    _zz_CtrlState_nextrndKey_610;
  wire       [1:0]    _zz_CtrlState_nextrndKey_611;
  wire       [1:0]    _zz_CtrlState_nextrndKey_612;
  wire                _zz_CtrlState_nextrndKey_613;
  reg        [1:0]    _zz_CtrlState_nextrndKey_614;
  wire       [1:0]    _zz_CtrlState_nextrndKey_615;
  reg        [1:0]    _zz_CtrlState_nextrndKey_616;
  wire                _zz_CtrlState_nextrndKey_617;
  reg        [1:0]    _zz_CtrlState_nextrndKey_618;
  wire                _zz_CtrlState_nextrndKey_619;
  reg        [1:0]    _zz_CtrlState_nextrndKey_620;
  wire       [7:0]    _zz_CtrlState_nextrndKey_621;
  reg        [7:0]    _zz_CtrlState_nextrndKey_622;
  wire                when_AES_CORE_l78;
  reg                 CtrlState_lastRound_regNext;
  (* ram_style = "distributed" *) reg [7:0] CtrlState_keyRcon [0:10];

  initial begin
    $readmemb("AES_CORE.v_toplevel_engine_CtrlState_keyRcon.bin",CtrlState_keyRcon);
  end
  assign _zz_CtrlState_keyRcon_port0 = CtrlState_keyRcon[_zz_CtrlState_nextrndKey_312];
  MyroundFunction rndFuc (
    .io_roundData (rndFuc_io_roundData[127:0]), //i
    .io_needMix   (rndFuc_io_needMix         ), //i
    .io_result    (rndFuc_io_result[127:0]   )  //o
  );
  assign CtrlState_lastRound = (CtrlState_rndCnt == 4'b1001);
  assign io_engine_cmd_fire = (io_engine_cmd_valid && io_engine_cmd_ready);
  always @(*) begin
    if(io_engine_cmd_fire) begin
      rndFuc_io_roundData = (io_engine_cmd_payload_block ^ CtrlState_currndKey);
    end else begin
      rndFuc_io_roundData = (CtrlState_dataBuf ^ CtrlState_currndKey);
    end
  end

  always @(*) begin
    if(io_engine_cmd_fire) begin
      rndFuc_io_needMix = (! CtrlState_lastRound);
    end else begin
      rndFuc_io_needMix = (! CtrlState_lastRound);
    end
  end

  always @(*) begin
    CtrlState_currndKey = 128'h0;
    if(io_engine_cmd_fire_1) begin
      CtrlState_currndKey = io_engine_cmd_payload_key;
    end else begin
      if(CtrlState_ongoing) begin
        CtrlState_currndKey = CtrlState_nextrndKey;
      end
    end
  end

  assign io_engine_cmd_fire_1 = (io_engine_cmd_valid && io_engine_cmd_ready);
  assign _zz_CtrlState_nextrndKey = {io_engine_cmd_payload_key[31 : 0],{io_engine_cmd_payload_key[63 : 32],{io_engine_cmd_payload_key[95 : 64],io_engine_cmd_payload_key[127 : 96]}}};
  assign _zz_CtrlState_nextrndKey_4 = _zz_CtrlState_nextrndKey[127 : 96];
  assign _zz_CtrlState_nextrndKey_5 = {_zz_CtrlState_nextrndKey_4[23 : 0],_zz_CtrlState_nextrndKey_4[31 : 24]};
  assign _zz_CtrlState_nextrndKey_7 = _zz_CtrlState_nextrndKey_5[7 : 0];
  always @(*) begin
    _zz_CtrlState_nextrndKey_10[7] = (((((_zz_CtrlState_nextrndKey_7[7] ^ _zz_CtrlState_nextrndKey_7[6]) ^ _zz_CtrlState_nextrndKey_7[5]) ^ _zz_CtrlState_nextrndKey_7[2]) ^ _zz_CtrlState_nextrndKey_7[1]) ^ _zz_CtrlState_nextrndKey_7[0]);
    _zz_CtrlState_nextrndKey_10[6] = (((_zz_CtrlState_nextrndKey_7[6] ^ _zz_CtrlState_nextrndKey_7[5]) ^ _zz_CtrlState_nextrndKey_7[4]) ^ _zz_CtrlState_nextrndKey_7[0]);
    _zz_CtrlState_nextrndKey_10[5] = (((_zz_CtrlState_nextrndKey_7[6] ^ _zz_CtrlState_nextrndKey_7[5]) ^ _zz_CtrlState_nextrndKey_7[1]) ^ _zz_CtrlState_nextrndKey_7[0]);
    _zz_CtrlState_nextrndKey_10[4] = (((_zz_CtrlState_nextrndKey_7[7] ^ _zz_CtrlState_nextrndKey_7[6]) ^ _zz_CtrlState_nextrndKey_7[5]) ^ _zz_CtrlState_nextrndKey_7[0]);
    _zz_CtrlState_nextrndKey_10[3] = ((((_zz_CtrlState_nextrndKey_7[7] ^ _zz_CtrlState_nextrndKey_7[4]) ^ _zz_CtrlState_nextrndKey_7[3]) ^ _zz_CtrlState_nextrndKey_7[1]) ^ _zz_CtrlState_nextrndKey_7[0]);
    _zz_CtrlState_nextrndKey_10[2] = _zz_CtrlState_nextrndKey_7[0];
    _zz_CtrlState_nextrndKey_10[1] = ((_zz_CtrlState_nextrndKey_7[6] ^ _zz_CtrlState_nextrndKey_7[5]) ^ _zz_CtrlState_nextrndKey_7[0]);
    _zz_CtrlState_nextrndKey_10[0] = ((((_zz_CtrlState_nextrndKey_7[6] ^ _zz_CtrlState_nextrndKey_7[3]) ^ _zz_CtrlState_nextrndKey_7[2]) ^ _zz_CtrlState_nextrndKey_7[1]) ^ _zz_CtrlState_nextrndKey_7[0]);
  end

  assign _zz_CtrlState_nextrndKey_9 = _zz_CtrlState_nextrndKey_10;
  assign _zz_CtrlState_nextrndKey_13 = _zz_CtrlState_nextrndKey_9[7 : 4];
  assign _zz_CtrlState_nextrndKey_14 = _zz_CtrlState_nextrndKey_9[3 : 0];
  assign _zz_CtrlState_nextrndKey_15 = (_zz_CtrlState_nextrndKey_13 ^ _zz_CtrlState_nextrndKey_14);
  always @(*) begin
    _zz_CtrlState_nextrndKey_16[3] = (_zz_CtrlState_nextrndKey_15[2] ^ _zz_CtrlState_nextrndKey_15[0]);
    _zz_CtrlState_nextrndKey_16[2] = (_zz_CtrlState_nextrndKey_15[3] ^ _zz_CtrlState_nextrndKey_15[1]);
    _zz_CtrlState_nextrndKey_16[1] = (_zz_CtrlState_nextrndKey_15[1] ^ _zz_CtrlState_nextrndKey_15[0]);
    _zz_CtrlState_nextrndKey_16[0] = _zz_CtrlState_nextrndKey_15[0];
  end

  assign _zz_CtrlState_nextrndKey_18 = _zz_CtrlState_nextrndKey_13[3 : 2];
  assign _zz_CtrlState_nextrndKey_19 = _zz_CtrlState_nextrndKey_13[1 : 0];
  assign _zz_CtrlState_nextrndKey_20 = _zz_CtrlState_nextrndKey_14[3 : 2];
  assign _zz_CtrlState_nextrndKey_21 = _zz_CtrlState_nextrndKey_14[1 : 0];
  assign _zz_CtrlState_nextrndKey_22 = (_zz_CtrlState_nextrndKey_18 ^ _zz_CtrlState_nextrndKey_19);
  assign _zz_CtrlState_nextrndKey_23 = (_zz_CtrlState_nextrndKey_20 ^ _zz_CtrlState_nextrndKey_21);
  assign _zz_CtrlState_nextrndKey_25 = ((_zz_CtrlState_nextrndKey_23[0] && _zz_CtrlState_nextrndKey_22[1]) ^ (_zz_CtrlState_nextrndKey_22[0] && _zz_CtrlState_nextrndKey_23[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_26[1] = ((_zz_CtrlState_nextrndKey_23[0] && _zz_CtrlState_nextrndKey_22[0]) ^ _zz_CtrlState_nextrndKey_25);
    _zz_CtrlState_nextrndKey_26[0] = ((_zz_CtrlState_nextrndKey_23[1] && _zz_CtrlState_nextrndKey_22[1]) ^ _zz_CtrlState_nextrndKey_25);
  end

  assign _zz_CtrlState_nextrndKey_24 = _zz_CtrlState_nextrndKey_26;
  always @(*) begin
    _zz_CtrlState_nextrndKey_28[1] = _zz_CtrlState_nextrndKey_24[0];
    _zz_CtrlState_nextrndKey_28[0] = (_zz_CtrlState_nextrndKey_24[0] ^ _zz_CtrlState_nextrndKey_24[1]);
  end

  assign _zz_CtrlState_nextrndKey_27 = _zz_CtrlState_nextrndKey_28;
  assign _zz_CtrlState_nextrndKey_29 = ((_zz_CtrlState_nextrndKey_20[0] && _zz_CtrlState_nextrndKey_18[1]) ^ (_zz_CtrlState_nextrndKey_18[0] && _zz_CtrlState_nextrndKey_20[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_30[1] = ((_zz_CtrlState_nextrndKey_20[0] && _zz_CtrlState_nextrndKey_18[0]) ^ _zz_CtrlState_nextrndKey_29);
    _zz_CtrlState_nextrndKey_30[0] = ((_zz_CtrlState_nextrndKey_20[1] && _zz_CtrlState_nextrndKey_18[1]) ^ _zz_CtrlState_nextrndKey_29);
  end

  assign _zz_CtrlState_nextrndKey_31 = ((_zz_CtrlState_nextrndKey_21[0] && _zz_CtrlState_nextrndKey_19[1]) ^ (_zz_CtrlState_nextrndKey_19[0] && _zz_CtrlState_nextrndKey_21[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_32[1] = ((_zz_CtrlState_nextrndKey_21[0] && _zz_CtrlState_nextrndKey_19[0]) ^ _zz_CtrlState_nextrndKey_31);
    _zz_CtrlState_nextrndKey_32[0] = ((_zz_CtrlState_nextrndKey_21[1] && _zz_CtrlState_nextrndKey_19[1]) ^ _zz_CtrlState_nextrndKey_31);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_17[3 : 2] = (_zz_CtrlState_nextrndKey_30 ^ _zz_CtrlState_nextrndKey_27);
    _zz_CtrlState_nextrndKey_17[1 : 0] = (_zz_CtrlState_nextrndKey_32 ^ _zz_CtrlState_nextrndKey_27);
  end

  assign _zz_CtrlState_nextrndKey_33 = (_zz_CtrlState_nextrndKey_16 ^ _zz_CtrlState_nextrndKey_17);
  assign _zz_CtrlState_nextrndKey_36 = _zz_CtrlState_nextrndKey_33[3 : 2];
  assign _zz_CtrlState_nextrndKey_37 = _zz_CtrlState_nextrndKey_33[1 : 0];
  assign _zz_CtrlState_nextrndKey_38 = (_zz_CtrlState_nextrndKey_36 ^ _zz_CtrlState_nextrndKey_37);
  always @(*) begin
    _zz_CtrlState_nextrndKey_39[1] = _zz_CtrlState_nextrndKey_38[1];
    _zz_CtrlState_nextrndKey_39[0] = (_zz_CtrlState_nextrndKey_38[0] ^ _zz_CtrlState_nextrndKey_38[1]);
  end

  assign _zz_CtrlState_nextrndKey_40 = ((_zz_CtrlState_nextrndKey_37[0] && _zz_CtrlState_nextrndKey_36[1]) ^ (_zz_CtrlState_nextrndKey_36[0] && _zz_CtrlState_nextrndKey_37[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_41[1] = ((_zz_CtrlState_nextrndKey_37[0] && _zz_CtrlState_nextrndKey_36[0]) ^ _zz_CtrlState_nextrndKey_40);
    _zz_CtrlState_nextrndKey_41[0] = ((_zz_CtrlState_nextrndKey_37[1] && _zz_CtrlState_nextrndKey_36[1]) ^ _zz_CtrlState_nextrndKey_40);
  end

  assign _zz_CtrlState_nextrndKey_42 = (_zz_CtrlState_nextrndKey_39 ^ _zz_CtrlState_nextrndKey_41);
  always @(*) begin
    _zz_CtrlState_nextrndKey_44[1] = _zz_CtrlState_nextrndKey_42[0];
    _zz_CtrlState_nextrndKey_44[0] = _zz_CtrlState_nextrndKey_42[1];
  end

  assign _zz_CtrlState_nextrndKey_43 = _zz_CtrlState_nextrndKey_44;
  assign _zz_CtrlState_nextrndKey_45 = ((_zz_CtrlState_nextrndKey_43[0] && _zz_CtrlState_nextrndKey_36[1]) ^ (_zz_CtrlState_nextrndKey_36[0] && _zz_CtrlState_nextrndKey_43[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_46[1] = ((_zz_CtrlState_nextrndKey_43[0] && _zz_CtrlState_nextrndKey_36[0]) ^ _zz_CtrlState_nextrndKey_45);
    _zz_CtrlState_nextrndKey_46[0] = ((_zz_CtrlState_nextrndKey_43[1] && _zz_CtrlState_nextrndKey_36[1]) ^ _zz_CtrlState_nextrndKey_45);
  end

  assign _zz_CtrlState_nextrndKey_47 = ((_zz_CtrlState_nextrndKey_43[0] && _zz_CtrlState_nextrndKey_37[1]) ^ (_zz_CtrlState_nextrndKey_37[0] && _zz_CtrlState_nextrndKey_43[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_48[1] = ((_zz_CtrlState_nextrndKey_43[0] && _zz_CtrlState_nextrndKey_37[0]) ^ _zz_CtrlState_nextrndKey_47);
    _zz_CtrlState_nextrndKey_48[0] = ((_zz_CtrlState_nextrndKey_43[1] && _zz_CtrlState_nextrndKey_37[1]) ^ _zz_CtrlState_nextrndKey_47);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_35[3 : 2] = _zz_CtrlState_nextrndKey_48;
    _zz_CtrlState_nextrndKey_35[1 : 0] = _zz_CtrlState_nextrndKey_46;
  end

  assign _zz_CtrlState_nextrndKey_34 = _zz_CtrlState_nextrndKey_35;
  assign _zz_CtrlState_nextrndKey_50 = _zz_CtrlState_nextrndKey_13[3 : 2];
  assign _zz_CtrlState_nextrndKey_51 = _zz_CtrlState_nextrndKey_13[1 : 0];
  assign _zz_CtrlState_nextrndKey_52 = _zz_CtrlState_nextrndKey_34[3 : 2];
  assign _zz_CtrlState_nextrndKey_53 = _zz_CtrlState_nextrndKey_34[1 : 0];
  assign _zz_CtrlState_nextrndKey_54 = (_zz_CtrlState_nextrndKey_50 ^ _zz_CtrlState_nextrndKey_51);
  assign _zz_CtrlState_nextrndKey_55 = (_zz_CtrlState_nextrndKey_52 ^ _zz_CtrlState_nextrndKey_53);
  assign _zz_CtrlState_nextrndKey_57 = ((_zz_CtrlState_nextrndKey_55[0] && _zz_CtrlState_nextrndKey_54[1]) ^ (_zz_CtrlState_nextrndKey_54[0] && _zz_CtrlState_nextrndKey_55[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_58[1] = ((_zz_CtrlState_nextrndKey_55[0] && _zz_CtrlState_nextrndKey_54[0]) ^ _zz_CtrlState_nextrndKey_57);
    _zz_CtrlState_nextrndKey_58[0] = ((_zz_CtrlState_nextrndKey_55[1] && _zz_CtrlState_nextrndKey_54[1]) ^ _zz_CtrlState_nextrndKey_57);
  end

  assign _zz_CtrlState_nextrndKey_56 = _zz_CtrlState_nextrndKey_58;
  always @(*) begin
    _zz_CtrlState_nextrndKey_60[1] = _zz_CtrlState_nextrndKey_56[0];
    _zz_CtrlState_nextrndKey_60[0] = (_zz_CtrlState_nextrndKey_56[0] ^ _zz_CtrlState_nextrndKey_56[1]);
  end

  assign _zz_CtrlState_nextrndKey_59 = _zz_CtrlState_nextrndKey_60;
  assign _zz_CtrlState_nextrndKey_61 = ((_zz_CtrlState_nextrndKey_52[0] && _zz_CtrlState_nextrndKey_50[1]) ^ (_zz_CtrlState_nextrndKey_50[0] && _zz_CtrlState_nextrndKey_52[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_62[1] = ((_zz_CtrlState_nextrndKey_52[0] && _zz_CtrlState_nextrndKey_50[0]) ^ _zz_CtrlState_nextrndKey_61);
    _zz_CtrlState_nextrndKey_62[0] = ((_zz_CtrlState_nextrndKey_52[1] && _zz_CtrlState_nextrndKey_50[1]) ^ _zz_CtrlState_nextrndKey_61);
  end

  assign _zz_CtrlState_nextrndKey_63 = ((_zz_CtrlState_nextrndKey_53[0] && _zz_CtrlState_nextrndKey_51[1]) ^ (_zz_CtrlState_nextrndKey_51[0] && _zz_CtrlState_nextrndKey_53[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_64[1] = ((_zz_CtrlState_nextrndKey_53[0] && _zz_CtrlState_nextrndKey_51[0]) ^ _zz_CtrlState_nextrndKey_63);
    _zz_CtrlState_nextrndKey_64[0] = ((_zz_CtrlState_nextrndKey_53[1] && _zz_CtrlState_nextrndKey_51[1]) ^ _zz_CtrlState_nextrndKey_63);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_49[3 : 2] = (_zz_CtrlState_nextrndKey_62 ^ _zz_CtrlState_nextrndKey_59);
    _zz_CtrlState_nextrndKey_49[1 : 0] = (_zz_CtrlState_nextrndKey_64 ^ _zz_CtrlState_nextrndKey_59);
  end

  assign _zz_CtrlState_nextrndKey_66 = _zz_CtrlState_nextrndKey_14[3 : 2];
  assign _zz_CtrlState_nextrndKey_67 = _zz_CtrlState_nextrndKey_14[1 : 0];
  assign _zz_CtrlState_nextrndKey_68 = _zz_CtrlState_nextrndKey_34[3 : 2];
  assign _zz_CtrlState_nextrndKey_69 = _zz_CtrlState_nextrndKey_34[1 : 0];
  assign _zz_CtrlState_nextrndKey_70 = (_zz_CtrlState_nextrndKey_66 ^ _zz_CtrlState_nextrndKey_67);
  assign _zz_CtrlState_nextrndKey_71 = (_zz_CtrlState_nextrndKey_68 ^ _zz_CtrlState_nextrndKey_69);
  assign _zz_CtrlState_nextrndKey_73 = ((_zz_CtrlState_nextrndKey_71[0] && _zz_CtrlState_nextrndKey_70[1]) ^ (_zz_CtrlState_nextrndKey_70[0] && _zz_CtrlState_nextrndKey_71[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_74[1] = ((_zz_CtrlState_nextrndKey_71[0] && _zz_CtrlState_nextrndKey_70[0]) ^ _zz_CtrlState_nextrndKey_73);
    _zz_CtrlState_nextrndKey_74[0] = ((_zz_CtrlState_nextrndKey_71[1] && _zz_CtrlState_nextrndKey_70[1]) ^ _zz_CtrlState_nextrndKey_73);
  end

  assign _zz_CtrlState_nextrndKey_72 = _zz_CtrlState_nextrndKey_74;
  always @(*) begin
    _zz_CtrlState_nextrndKey_76[1] = _zz_CtrlState_nextrndKey_72[0];
    _zz_CtrlState_nextrndKey_76[0] = (_zz_CtrlState_nextrndKey_72[0] ^ _zz_CtrlState_nextrndKey_72[1]);
  end

  assign _zz_CtrlState_nextrndKey_75 = _zz_CtrlState_nextrndKey_76;
  assign _zz_CtrlState_nextrndKey_77 = ((_zz_CtrlState_nextrndKey_68[0] && _zz_CtrlState_nextrndKey_66[1]) ^ (_zz_CtrlState_nextrndKey_66[0] && _zz_CtrlState_nextrndKey_68[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_78[1] = ((_zz_CtrlState_nextrndKey_68[0] && _zz_CtrlState_nextrndKey_66[0]) ^ _zz_CtrlState_nextrndKey_77);
    _zz_CtrlState_nextrndKey_78[0] = ((_zz_CtrlState_nextrndKey_68[1] && _zz_CtrlState_nextrndKey_66[1]) ^ _zz_CtrlState_nextrndKey_77);
  end

  assign _zz_CtrlState_nextrndKey_79 = ((_zz_CtrlState_nextrndKey_69[0] && _zz_CtrlState_nextrndKey_67[1]) ^ (_zz_CtrlState_nextrndKey_67[0] && _zz_CtrlState_nextrndKey_69[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_80[1] = ((_zz_CtrlState_nextrndKey_69[0] && _zz_CtrlState_nextrndKey_67[0]) ^ _zz_CtrlState_nextrndKey_79);
    _zz_CtrlState_nextrndKey_80[0] = ((_zz_CtrlState_nextrndKey_69[1] && _zz_CtrlState_nextrndKey_67[1]) ^ _zz_CtrlState_nextrndKey_79);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_65[3 : 2] = (_zz_CtrlState_nextrndKey_78 ^ _zz_CtrlState_nextrndKey_75);
    _zz_CtrlState_nextrndKey_65[1 : 0] = (_zz_CtrlState_nextrndKey_80 ^ _zz_CtrlState_nextrndKey_75);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_12[7 : 4] = _zz_CtrlState_nextrndKey_65;
    _zz_CtrlState_nextrndKey_12[3 : 0] = _zz_CtrlState_nextrndKey_49;
  end

  assign _zz_CtrlState_nextrndKey_11 = _zz_CtrlState_nextrndKey_12;
  always @(*) begin
    _zz_CtrlState_nextrndKey_82[7] = (_zz_CtrlState_nextrndKey_11[5] ^ _zz_CtrlState_nextrndKey_11[3]);
    _zz_CtrlState_nextrndKey_82[6] = (_zz_CtrlState_nextrndKey_11[7] ^ _zz_CtrlState_nextrndKey_11[3]);
    _zz_CtrlState_nextrndKey_82[5] = (_zz_CtrlState_nextrndKey_11[6] ^ _zz_CtrlState_nextrndKey_11[0]);
    _zz_CtrlState_nextrndKey_82[4] = ((_zz_CtrlState_nextrndKey_11[7] ^ _zz_CtrlState_nextrndKey_11[5]) ^ _zz_CtrlState_nextrndKey_11[3]);
    _zz_CtrlState_nextrndKey_82[3] = ((((_zz_CtrlState_nextrndKey_11[7] ^ _zz_CtrlState_nextrndKey_11[6]) ^ _zz_CtrlState_nextrndKey_11[5]) ^ _zz_CtrlState_nextrndKey_11[4]) ^ _zz_CtrlState_nextrndKey_11[3]);
    _zz_CtrlState_nextrndKey_82[2] = ((((_zz_CtrlState_nextrndKey_11[6] ^ _zz_CtrlState_nextrndKey_11[5]) ^ _zz_CtrlState_nextrndKey_11[3]) ^ _zz_CtrlState_nextrndKey_11[2]) ^ _zz_CtrlState_nextrndKey_11[0]);
    _zz_CtrlState_nextrndKey_82[1] = ((_zz_CtrlState_nextrndKey_11[5] ^ _zz_CtrlState_nextrndKey_11[4]) ^ _zz_CtrlState_nextrndKey_11[1]);
    _zz_CtrlState_nextrndKey_82[0] = ((_zz_CtrlState_nextrndKey_11[6] ^ _zz_CtrlState_nextrndKey_11[4]) ^ _zz_CtrlState_nextrndKey_11[1]);
  end

  assign _zz_CtrlState_nextrndKey_81 = _zz_CtrlState_nextrndKey_82;
  always @(*) begin
    _zz_CtrlState_nextrndKey_8[7] = _zz_CtrlState_nextrndKey_81[7];
    _zz_CtrlState_nextrndKey_8[6] = (! _zz_CtrlState_nextrndKey_81[6]);
    _zz_CtrlState_nextrndKey_8[5] = (! _zz_CtrlState_nextrndKey_81[5]);
    _zz_CtrlState_nextrndKey_8[4] = _zz_CtrlState_nextrndKey_81[4];
    _zz_CtrlState_nextrndKey_8[3] = _zz_CtrlState_nextrndKey_81[3];
    _zz_CtrlState_nextrndKey_8[2] = _zz_CtrlState_nextrndKey_81[2];
    _zz_CtrlState_nextrndKey_8[1] = (! _zz_CtrlState_nextrndKey_81[1]);
    _zz_CtrlState_nextrndKey_8[0] = (! _zz_CtrlState_nextrndKey_81[0]);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_6[7 : 0] = _zz_CtrlState_nextrndKey_8;
    _zz_CtrlState_nextrndKey_6[15 : 8] = _zz_CtrlState_nextrndKey_84;
    _zz_CtrlState_nextrndKey_6[23 : 16] = _zz_CtrlState_nextrndKey_160;
    _zz_CtrlState_nextrndKey_6[31 : 24] = _zz_CtrlState_nextrndKey_236;
  end

  assign _zz_CtrlState_nextrndKey_83 = _zz_CtrlState_nextrndKey_5[15 : 8];
  always @(*) begin
    _zz_CtrlState_nextrndKey_86[7] = (((((_zz_CtrlState_nextrndKey_83[7] ^ _zz_CtrlState_nextrndKey_83[6]) ^ _zz_CtrlState_nextrndKey_83[5]) ^ _zz_CtrlState_nextrndKey_83[2]) ^ _zz_CtrlState_nextrndKey_83[1]) ^ _zz_CtrlState_nextrndKey_83[0]);
    _zz_CtrlState_nextrndKey_86[6] = (((_zz_CtrlState_nextrndKey_83[6] ^ _zz_CtrlState_nextrndKey_83[5]) ^ _zz_CtrlState_nextrndKey_83[4]) ^ _zz_CtrlState_nextrndKey_83[0]);
    _zz_CtrlState_nextrndKey_86[5] = (((_zz_CtrlState_nextrndKey_83[6] ^ _zz_CtrlState_nextrndKey_83[5]) ^ _zz_CtrlState_nextrndKey_83[1]) ^ _zz_CtrlState_nextrndKey_83[0]);
    _zz_CtrlState_nextrndKey_86[4] = (((_zz_CtrlState_nextrndKey_83[7] ^ _zz_CtrlState_nextrndKey_83[6]) ^ _zz_CtrlState_nextrndKey_83[5]) ^ _zz_CtrlState_nextrndKey_83[0]);
    _zz_CtrlState_nextrndKey_86[3] = ((((_zz_CtrlState_nextrndKey_83[7] ^ _zz_CtrlState_nextrndKey_83[4]) ^ _zz_CtrlState_nextrndKey_83[3]) ^ _zz_CtrlState_nextrndKey_83[1]) ^ _zz_CtrlState_nextrndKey_83[0]);
    _zz_CtrlState_nextrndKey_86[2] = _zz_CtrlState_nextrndKey_83[0];
    _zz_CtrlState_nextrndKey_86[1] = ((_zz_CtrlState_nextrndKey_83[6] ^ _zz_CtrlState_nextrndKey_83[5]) ^ _zz_CtrlState_nextrndKey_83[0]);
    _zz_CtrlState_nextrndKey_86[0] = ((((_zz_CtrlState_nextrndKey_83[6] ^ _zz_CtrlState_nextrndKey_83[3]) ^ _zz_CtrlState_nextrndKey_83[2]) ^ _zz_CtrlState_nextrndKey_83[1]) ^ _zz_CtrlState_nextrndKey_83[0]);
  end

  assign _zz_CtrlState_nextrndKey_85 = _zz_CtrlState_nextrndKey_86;
  assign _zz_CtrlState_nextrndKey_89 = _zz_CtrlState_nextrndKey_85[7 : 4];
  assign _zz_CtrlState_nextrndKey_90 = _zz_CtrlState_nextrndKey_85[3 : 0];
  assign _zz_CtrlState_nextrndKey_91 = (_zz_CtrlState_nextrndKey_89 ^ _zz_CtrlState_nextrndKey_90);
  always @(*) begin
    _zz_CtrlState_nextrndKey_92[3] = (_zz_CtrlState_nextrndKey_91[2] ^ _zz_CtrlState_nextrndKey_91[0]);
    _zz_CtrlState_nextrndKey_92[2] = (_zz_CtrlState_nextrndKey_91[3] ^ _zz_CtrlState_nextrndKey_91[1]);
    _zz_CtrlState_nextrndKey_92[1] = (_zz_CtrlState_nextrndKey_91[1] ^ _zz_CtrlState_nextrndKey_91[0]);
    _zz_CtrlState_nextrndKey_92[0] = _zz_CtrlState_nextrndKey_91[0];
  end

  assign _zz_CtrlState_nextrndKey_94 = _zz_CtrlState_nextrndKey_89[3 : 2];
  assign _zz_CtrlState_nextrndKey_95 = _zz_CtrlState_nextrndKey_89[1 : 0];
  assign _zz_CtrlState_nextrndKey_96 = _zz_CtrlState_nextrndKey_90[3 : 2];
  assign _zz_CtrlState_nextrndKey_97 = _zz_CtrlState_nextrndKey_90[1 : 0];
  assign _zz_CtrlState_nextrndKey_98 = (_zz_CtrlState_nextrndKey_94 ^ _zz_CtrlState_nextrndKey_95);
  assign _zz_CtrlState_nextrndKey_99 = (_zz_CtrlState_nextrndKey_96 ^ _zz_CtrlState_nextrndKey_97);
  assign _zz_CtrlState_nextrndKey_101 = ((_zz_CtrlState_nextrndKey_99[0] && _zz_CtrlState_nextrndKey_98[1]) ^ (_zz_CtrlState_nextrndKey_98[0] && _zz_CtrlState_nextrndKey_99[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_102[1] = ((_zz_CtrlState_nextrndKey_99[0] && _zz_CtrlState_nextrndKey_98[0]) ^ _zz_CtrlState_nextrndKey_101);
    _zz_CtrlState_nextrndKey_102[0] = ((_zz_CtrlState_nextrndKey_99[1] && _zz_CtrlState_nextrndKey_98[1]) ^ _zz_CtrlState_nextrndKey_101);
  end

  assign _zz_CtrlState_nextrndKey_100 = _zz_CtrlState_nextrndKey_102;
  always @(*) begin
    _zz_CtrlState_nextrndKey_104[1] = _zz_CtrlState_nextrndKey_100[0];
    _zz_CtrlState_nextrndKey_104[0] = (_zz_CtrlState_nextrndKey_100[0] ^ _zz_CtrlState_nextrndKey_100[1]);
  end

  assign _zz_CtrlState_nextrndKey_103 = _zz_CtrlState_nextrndKey_104;
  assign _zz_CtrlState_nextrndKey_105 = ((_zz_CtrlState_nextrndKey_96[0] && _zz_CtrlState_nextrndKey_94[1]) ^ (_zz_CtrlState_nextrndKey_94[0] && _zz_CtrlState_nextrndKey_96[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_106[1] = ((_zz_CtrlState_nextrndKey_96[0] && _zz_CtrlState_nextrndKey_94[0]) ^ _zz_CtrlState_nextrndKey_105);
    _zz_CtrlState_nextrndKey_106[0] = ((_zz_CtrlState_nextrndKey_96[1] && _zz_CtrlState_nextrndKey_94[1]) ^ _zz_CtrlState_nextrndKey_105);
  end

  assign _zz_CtrlState_nextrndKey_107 = ((_zz_CtrlState_nextrndKey_97[0] && _zz_CtrlState_nextrndKey_95[1]) ^ (_zz_CtrlState_nextrndKey_95[0] && _zz_CtrlState_nextrndKey_97[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_108[1] = ((_zz_CtrlState_nextrndKey_97[0] && _zz_CtrlState_nextrndKey_95[0]) ^ _zz_CtrlState_nextrndKey_107);
    _zz_CtrlState_nextrndKey_108[0] = ((_zz_CtrlState_nextrndKey_97[1] && _zz_CtrlState_nextrndKey_95[1]) ^ _zz_CtrlState_nextrndKey_107);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_93[3 : 2] = (_zz_CtrlState_nextrndKey_106 ^ _zz_CtrlState_nextrndKey_103);
    _zz_CtrlState_nextrndKey_93[1 : 0] = (_zz_CtrlState_nextrndKey_108 ^ _zz_CtrlState_nextrndKey_103);
  end

  assign _zz_CtrlState_nextrndKey_109 = (_zz_CtrlState_nextrndKey_92 ^ _zz_CtrlState_nextrndKey_93);
  assign _zz_CtrlState_nextrndKey_112 = _zz_CtrlState_nextrndKey_109[3 : 2];
  assign _zz_CtrlState_nextrndKey_113 = _zz_CtrlState_nextrndKey_109[1 : 0];
  assign _zz_CtrlState_nextrndKey_114 = (_zz_CtrlState_nextrndKey_112 ^ _zz_CtrlState_nextrndKey_113);
  always @(*) begin
    _zz_CtrlState_nextrndKey_115[1] = _zz_CtrlState_nextrndKey_114[1];
    _zz_CtrlState_nextrndKey_115[0] = (_zz_CtrlState_nextrndKey_114[0] ^ _zz_CtrlState_nextrndKey_114[1]);
  end

  assign _zz_CtrlState_nextrndKey_116 = ((_zz_CtrlState_nextrndKey_113[0] && _zz_CtrlState_nextrndKey_112[1]) ^ (_zz_CtrlState_nextrndKey_112[0] && _zz_CtrlState_nextrndKey_113[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_117[1] = ((_zz_CtrlState_nextrndKey_113[0] && _zz_CtrlState_nextrndKey_112[0]) ^ _zz_CtrlState_nextrndKey_116);
    _zz_CtrlState_nextrndKey_117[0] = ((_zz_CtrlState_nextrndKey_113[1] && _zz_CtrlState_nextrndKey_112[1]) ^ _zz_CtrlState_nextrndKey_116);
  end

  assign _zz_CtrlState_nextrndKey_118 = (_zz_CtrlState_nextrndKey_115 ^ _zz_CtrlState_nextrndKey_117);
  always @(*) begin
    _zz_CtrlState_nextrndKey_120[1] = _zz_CtrlState_nextrndKey_118[0];
    _zz_CtrlState_nextrndKey_120[0] = _zz_CtrlState_nextrndKey_118[1];
  end

  assign _zz_CtrlState_nextrndKey_119 = _zz_CtrlState_nextrndKey_120;
  assign _zz_CtrlState_nextrndKey_121 = ((_zz_CtrlState_nextrndKey_119[0] && _zz_CtrlState_nextrndKey_112[1]) ^ (_zz_CtrlState_nextrndKey_112[0] && _zz_CtrlState_nextrndKey_119[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_122[1] = ((_zz_CtrlState_nextrndKey_119[0] && _zz_CtrlState_nextrndKey_112[0]) ^ _zz_CtrlState_nextrndKey_121);
    _zz_CtrlState_nextrndKey_122[0] = ((_zz_CtrlState_nextrndKey_119[1] && _zz_CtrlState_nextrndKey_112[1]) ^ _zz_CtrlState_nextrndKey_121);
  end

  assign _zz_CtrlState_nextrndKey_123 = ((_zz_CtrlState_nextrndKey_119[0] && _zz_CtrlState_nextrndKey_113[1]) ^ (_zz_CtrlState_nextrndKey_113[0] && _zz_CtrlState_nextrndKey_119[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_124[1] = ((_zz_CtrlState_nextrndKey_119[0] && _zz_CtrlState_nextrndKey_113[0]) ^ _zz_CtrlState_nextrndKey_123);
    _zz_CtrlState_nextrndKey_124[0] = ((_zz_CtrlState_nextrndKey_119[1] && _zz_CtrlState_nextrndKey_113[1]) ^ _zz_CtrlState_nextrndKey_123);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_111[3 : 2] = _zz_CtrlState_nextrndKey_124;
    _zz_CtrlState_nextrndKey_111[1 : 0] = _zz_CtrlState_nextrndKey_122;
  end

  assign _zz_CtrlState_nextrndKey_110 = _zz_CtrlState_nextrndKey_111;
  assign _zz_CtrlState_nextrndKey_126 = _zz_CtrlState_nextrndKey_89[3 : 2];
  assign _zz_CtrlState_nextrndKey_127 = _zz_CtrlState_nextrndKey_89[1 : 0];
  assign _zz_CtrlState_nextrndKey_128 = _zz_CtrlState_nextrndKey_110[3 : 2];
  assign _zz_CtrlState_nextrndKey_129 = _zz_CtrlState_nextrndKey_110[1 : 0];
  assign _zz_CtrlState_nextrndKey_130 = (_zz_CtrlState_nextrndKey_126 ^ _zz_CtrlState_nextrndKey_127);
  assign _zz_CtrlState_nextrndKey_131 = (_zz_CtrlState_nextrndKey_128 ^ _zz_CtrlState_nextrndKey_129);
  assign _zz_CtrlState_nextrndKey_133 = ((_zz_CtrlState_nextrndKey_131[0] && _zz_CtrlState_nextrndKey_130[1]) ^ (_zz_CtrlState_nextrndKey_130[0] && _zz_CtrlState_nextrndKey_131[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_134[1] = ((_zz_CtrlState_nextrndKey_131[0] && _zz_CtrlState_nextrndKey_130[0]) ^ _zz_CtrlState_nextrndKey_133);
    _zz_CtrlState_nextrndKey_134[0] = ((_zz_CtrlState_nextrndKey_131[1] && _zz_CtrlState_nextrndKey_130[1]) ^ _zz_CtrlState_nextrndKey_133);
  end

  assign _zz_CtrlState_nextrndKey_132 = _zz_CtrlState_nextrndKey_134;
  always @(*) begin
    _zz_CtrlState_nextrndKey_136[1] = _zz_CtrlState_nextrndKey_132[0];
    _zz_CtrlState_nextrndKey_136[0] = (_zz_CtrlState_nextrndKey_132[0] ^ _zz_CtrlState_nextrndKey_132[1]);
  end

  assign _zz_CtrlState_nextrndKey_135 = _zz_CtrlState_nextrndKey_136;
  assign _zz_CtrlState_nextrndKey_137 = ((_zz_CtrlState_nextrndKey_128[0] && _zz_CtrlState_nextrndKey_126[1]) ^ (_zz_CtrlState_nextrndKey_126[0] && _zz_CtrlState_nextrndKey_128[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_138[1] = ((_zz_CtrlState_nextrndKey_128[0] && _zz_CtrlState_nextrndKey_126[0]) ^ _zz_CtrlState_nextrndKey_137);
    _zz_CtrlState_nextrndKey_138[0] = ((_zz_CtrlState_nextrndKey_128[1] && _zz_CtrlState_nextrndKey_126[1]) ^ _zz_CtrlState_nextrndKey_137);
  end

  assign _zz_CtrlState_nextrndKey_139 = ((_zz_CtrlState_nextrndKey_129[0] && _zz_CtrlState_nextrndKey_127[1]) ^ (_zz_CtrlState_nextrndKey_127[0] && _zz_CtrlState_nextrndKey_129[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_140[1] = ((_zz_CtrlState_nextrndKey_129[0] && _zz_CtrlState_nextrndKey_127[0]) ^ _zz_CtrlState_nextrndKey_139);
    _zz_CtrlState_nextrndKey_140[0] = ((_zz_CtrlState_nextrndKey_129[1] && _zz_CtrlState_nextrndKey_127[1]) ^ _zz_CtrlState_nextrndKey_139);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_125[3 : 2] = (_zz_CtrlState_nextrndKey_138 ^ _zz_CtrlState_nextrndKey_135);
    _zz_CtrlState_nextrndKey_125[1 : 0] = (_zz_CtrlState_nextrndKey_140 ^ _zz_CtrlState_nextrndKey_135);
  end

  assign _zz_CtrlState_nextrndKey_142 = _zz_CtrlState_nextrndKey_90[3 : 2];
  assign _zz_CtrlState_nextrndKey_143 = _zz_CtrlState_nextrndKey_90[1 : 0];
  assign _zz_CtrlState_nextrndKey_144 = _zz_CtrlState_nextrndKey_110[3 : 2];
  assign _zz_CtrlState_nextrndKey_145 = _zz_CtrlState_nextrndKey_110[1 : 0];
  assign _zz_CtrlState_nextrndKey_146 = (_zz_CtrlState_nextrndKey_142 ^ _zz_CtrlState_nextrndKey_143);
  assign _zz_CtrlState_nextrndKey_147 = (_zz_CtrlState_nextrndKey_144 ^ _zz_CtrlState_nextrndKey_145);
  assign _zz_CtrlState_nextrndKey_149 = ((_zz_CtrlState_nextrndKey_147[0] && _zz_CtrlState_nextrndKey_146[1]) ^ (_zz_CtrlState_nextrndKey_146[0] && _zz_CtrlState_nextrndKey_147[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_150[1] = ((_zz_CtrlState_nextrndKey_147[0] && _zz_CtrlState_nextrndKey_146[0]) ^ _zz_CtrlState_nextrndKey_149);
    _zz_CtrlState_nextrndKey_150[0] = ((_zz_CtrlState_nextrndKey_147[1] && _zz_CtrlState_nextrndKey_146[1]) ^ _zz_CtrlState_nextrndKey_149);
  end

  assign _zz_CtrlState_nextrndKey_148 = _zz_CtrlState_nextrndKey_150;
  always @(*) begin
    _zz_CtrlState_nextrndKey_152[1] = _zz_CtrlState_nextrndKey_148[0];
    _zz_CtrlState_nextrndKey_152[0] = (_zz_CtrlState_nextrndKey_148[0] ^ _zz_CtrlState_nextrndKey_148[1]);
  end

  assign _zz_CtrlState_nextrndKey_151 = _zz_CtrlState_nextrndKey_152;
  assign _zz_CtrlState_nextrndKey_153 = ((_zz_CtrlState_nextrndKey_144[0] && _zz_CtrlState_nextrndKey_142[1]) ^ (_zz_CtrlState_nextrndKey_142[0] && _zz_CtrlState_nextrndKey_144[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_154[1] = ((_zz_CtrlState_nextrndKey_144[0] && _zz_CtrlState_nextrndKey_142[0]) ^ _zz_CtrlState_nextrndKey_153);
    _zz_CtrlState_nextrndKey_154[0] = ((_zz_CtrlState_nextrndKey_144[1] && _zz_CtrlState_nextrndKey_142[1]) ^ _zz_CtrlState_nextrndKey_153);
  end

  assign _zz_CtrlState_nextrndKey_155 = ((_zz_CtrlState_nextrndKey_145[0] && _zz_CtrlState_nextrndKey_143[1]) ^ (_zz_CtrlState_nextrndKey_143[0] && _zz_CtrlState_nextrndKey_145[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_156[1] = ((_zz_CtrlState_nextrndKey_145[0] && _zz_CtrlState_nextrndKey_143[0]) ^ _zz_CtrlState_nextrndKey_155);
    _zz_CtrlState_nextrndKey_156[0] = ((_zz_CtrlState_nextrndKey_145[1] && _zz_CtrlState_nextrndKey_143[1]) ^ _zz_CtrlState_nextrndKey_155);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_141[3 : 2] = (_zz_CtrlState_nextrndKey_154 ^ _zz_CtrlState_nextrndKey_151);
    _zz_CtrlState_nextrndKey_141[1 : 0] = (_zz_CtrlState_nextrndKey_156 ^ _zz_CtrlState_nextrndKey_151);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_88[7 : 4] = _zz_CtrlState_nextrndKey_141;
    _zz_CtrlState_nextrndKey_88[3 : 0] = _zz_CtrlState_nextrndKey_125;
  end

  assign _zz_CtrlState_nextrndKey_87 = _zz_CtrlState_nextrndKey_88;
  always @(*) begin
    _zz_CtrlState_nextrndKey_158[7] = (_zz_CtrlState_nextrndKey_87[5] ^ _zz_CtrlState_nextrndKey_87[3]);
    _zz_CtrlState_nextrndKey_158[6] = (_zz_CtrlState_nextrndKey_87[7] ^ _zz_CtrlState_nextrndKey_87[3]);
    _zz_CtrlState_nextrndKey_158[5] = (_zz_CtrlState_nextrndKey_87[6] ^ _zz_CtrlState_nextrndKey_87[0]);
    _zz_CtrlState_nextrndKey_158[4] = ((_zz_CtrlState_nextrndKey_87[7] ^ _zz_CtrlState_nextrndKey_87[5]) ^ _zz_CtrlState_nextrndKey_87[3]);
    _zz_CtrlState_nextrndKey_158[3] = ((((_zz_CtrlState_nextrndKey_87[7] ^ _zz_CtrlState_nextrndKey_87[6]) ^ _zz_CtrlState_nextrndKey_87[5]) ^ _zz_CtrlState_nextrndKey_87[4]) ^ _zz_CtrlState_nextrndKey_87[3]);
    _zz_CtrlState_nextrndKey_158[2] = ((((_zz_CtrlState_nextrndKey_87[6] ^ _zz_CtrlState_nextrndKey_87[5]) ^ _zz_CtrlState_nextrndKey_87[3]) ^ _zz_CtrlState_nextrndKey_87[2]) ^ _zz_CtrlState_nextrndKey_87[0]);
    _zz_CtrlState_nextrndKey_158[1] = ((_zz_CtrlState_nextrndKey_87[5] ^ _zz_CtrlState_nextrndKey_87[4]) ^ _zz_CtrlState_nextrndKey_87[1]);
    _zz_CtrlState_nextrndKey_158[0] = ((_zz_CtrlState_nextrndKey_87[6] ^ _zz_CtrlState_nextrndKey_87[4]) ^ _zz_CtrlState_nextrndKey_87[1]);
  end

  assign _zz_CtrlState_nextrndKey_157 = _zz_CtrlState_nextrndKey_158;
  always @(*) begin
    _zz_CtrlState_nextrndKey_84[7] = _zz_CtrlState_nextrndKey_157[7];
    _zz_CtrlState_nextrndKey_84[6] = (! _zz_CtrlState_nextrndKey_157[6]);
    _zz_CtrlState_nextrndKey_84[5] = (! _zz_CtrlState_nextrndKey_157[5]);
    _zz_CtrlState_nextrndKey_84[4] = _zz_CtrlState_nextrndKey_157[4];
    _zz_CtrlState_nextrndKey_84[3] = _zz_CtrlState_nextrndKey_157[3];
    _zz_CtrlState_nextrndKey_84[2] = _zz_CtrlState_nextrndKey_157[2];
    _zz_CtrlState_nextrndKey_84[1] = (! _zz_CtrlState_nextrndKey_157[1]);
    _zz_CtrlState_nextrndKey_84[0] = (! _zz_CtrlState_nextrndKey_157[0]);
  end

  assign _zz_CtrlState_nextrndKey_159 = _zz_CtrlState_nextrndKey_5[23 : 16];
  always @(*) begin
    _zz_CtrlState_nextrndKey_162[7] = (((((_zz_CtrlState_nextrndKey_159[7] ^ _zz_CtrlState_nextrndKey_159[6]) ^ _zz_CtrlState_nextrndKey_159[5]) ^ _zz_CtrlState_nextrndKey_159[2]) ^ _zz_CtrlState_nextrndKey_159[1]) ^ _zz_CtrlState_nextrndKey_159[0]);
    _zz_CtrlState_nextrndKey_162[6] = (((_zz_CtrlState_nextrndKey_159[6] ^ _zz_CtrlState_nextrndKey_159[5]) ^ _zz_CtrlState_nextrndKey_159[4]) ^ _zz_CtrlState_nextrndKey_159[0]);
    _zz_CtrlState_nextrndKey_162[5] = (((_zz_CtrlState_nextrndKey_159[6] ^ _zz_CtrlState_nextrndKey_159[5]) ^ _zz_CtrlState_nextrndKey_159[1]) ^ _zz_CtrlState_nextrndKey_159[0]);
    _zz_CtrlState_nextrndKey_162[4] = (((_zz_CtrlState_nextrndKey_159[7] ^ _zz_CtrlState_nextrndKey_159[6]) ^ _zz_CtrlState_nextrndKey_159[5]) ^ _zz_CtrlState_nextrndKey_159[0]);
    _zz_CtrlState_nextrndKey_162[3] = ((((_zz_CtrlState_nextrndKey_159[7] ^ _zz_CtrlState_nextrndKey_159[4]) ^ _zz_CtrlState_nextrndKey_159[3]) ^ _zz_CtrlState_nextrndKey_159[1]) ^ _zz_CtrlState_nextrndKey_159[0]);
    _zz_CtrlState_nextrndKey_162[2] = _zz_CtrlState_nextrndKey_159[0];
    _zz_CtrlState_nextrndKey_162[1] = ((_zz_CtrlState_nextrndKey_159[6] ^ _zz_CtrlState_nextrndKey_159[5]) ^ _zz_CtrlState_nextrndKey_159[0]);
    _zz_CtrlState_nextrndKey_162[0] = ((((_zz_CtrlState_nextrndKey_159[6] ^ _zz_CtrlState_nextrndKey_159[3]) ^ _zz_CtrlState_nextrndKey_159[2]) ^ _zz_CtrlState_nextrndKey_159[1]) ^ _zz_CtrlState_nextrndKey_159[0]);
  end

  assign _zz_CtrlState_nextrndKey_161 = _zz_CtrlState_nextrndKey_162;
  assign _zz_CtrlState_nextrndKey_165 = _zz_CtrlState_nextrndKey_161[7 : 4];
  assign _zz_CtrlState_nextrndKey_166 = _zz_CtrlState_nextrndKey_161[3 : 0];
  assign _zz_CtrlState_nextrndKey_167 = (_zz_CtrlState_nextrndKey_165 ^ _zz_CtrlState_nextrndKey_166);
  always @(*) begin
    _zz_CtrlState_nextrndKey_168[3] = (_zz_CtrlState_nextrndKey_167[2] ^ _zz_CtrlState_nextrndKey_167[0]);
    _zz_CtrlState_nextrndKey_168[2] = (_zz_CtrlState_nextrndKey_167[3] ^ _zz_CtrlState_nextrndKey_167[1]);
    _zz_CtrlState_nextrndKey_168[1] = (_zz_CtrlState_nextrndKey_167[1] ^ _zz_CtrlState_nextrndKey_167[0]);
    _zz_CtrlState_nextrndKey_168[0] = _zz_CtrlState_nextrndKey_167[0];
  end

  assign _zz_CtrlState_nextrndKey_170 = _zz_CtrlState_nextrndKey_165[3 : 2];
  assign _zz_CtrlState_nextrndKey_171 = _zz_CtrlState_nextrndKey_165[1 : 0];
  assign _zz_CtrlState_nextrndKey_172 = _zz_CtrlState_nextrndKey_166[3 : 2];
  assign _zz_CtrlState_nextrndKey_173 = _zz_CtrlState_nextrndKey_166[1 : 0];
  assign _zz_CtrlState_nextrndKey_174 = (_zz_CtrlState_nextrndKey_170 ^ _zz_CtrlState_nextrndKey_171);
  assign _zz_CtrlState_nextrndKey_175 = (_zz_CtrlState_nextrndKey_172 ^ _zz_CtrlState_nextrndKey_173);
  assign _zz_CtrlState_nextrndKey_177 = ((_zz_CtrlState_nextrndKey_175[0] && _zz_CtrlState_nextrndKey_174[1]) ^ (_zz_CtrlState_nextrndKey_174[0] && _zz_CtrlState_nextrndKey_175[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_178[1] = ((_zz_CtrlState_nextrndKey_175[0] && _zz_CtrlState_nextrndKey_174[0]) ^ _zz_CtrlState_nextrndKey_177);
    _zz_CtrlState_nextrndKey_178[0] = ((_zz_CtrlState_nextrndKey_175[1] && _zz_CtrlState_nextrndKey_174[1]) ^ _zz_CtrlState_nextrndKey_177);
  end

  assign _zz_CtrlState_nextrndKey_176 = _zz_CtrlState_nextrndKey_178;
  always @(*) begin
    _zz_CtrlState_nextrndKey_180[1] = _zz_CtrlState_nextrndKey_176[0];
    _zz_CtrlState_nextrndKey_180[0] = (_zz_CtrlState_nextrndKey_176[0] ^ _zz_CtrlState_nextrndKey_176[1]);
  end

  assign _zz_CtrlState_nextrndKey_179 = _zz_CtrlState_nextrndKey_180;
  assign _zz_CtrlState_nextrndKey_181 = ((_zz_CtrlState_nextrndKey_172[0] && _zz_CtrlState_nextrndKey_170[1]) ^ (_zz_CtrlState_nextrndKey_170[0] && _zz_CtrlState_nextrndKey_172[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_182[1] = ((_zz_CtrlState_nextrndKey_172[0] && _zz_CtrlState_nextrndKey_170[0]) ^ _zz_CtrlState_nextrndKey_181);
    _zz_CtrlState_nextrndKey_182[0] = ((_zz_CtrlState_nextrndKey_172[1] && _zz_CtrlState_nextrndKey_170[1]) ^ _zz_CtrlState_nextrndKey_181);
  end

  assign _zz_CtrlState_nextrndKey_183 = ((_zz_CtrlState_nextrndKey_173[0] && _zz_CtrlState_nextrndKey_171[1]) ^ (_zz_CtrlState_nextrndKey_171[0] && _zz_CtrlState_nextrndKey_173[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_184[1] = ((_zz_CtrlState_nextrndKey_173[0] && _zz_CtrlState_nextrndKey_171[0]) ^ _zz_CtrlState_nextrndKey_183);
    _zz_CtrlState_nextrndKey_184[0] = ((_zz_CtrlState_nextrndKey_173[1] && _zz_CtrlState_nextrndKey_171[1]) ^ _zz_CtrlState_nextrndKey_183);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_169[3 : 2] = (_zz_CtrlState_nextrndKey_182 ^ _zz_CtrlState_nextrndKey_179);
    _zz_CtrlState_nextrndKey_169[1 : 0] = (_zz_CtrlState_nextrndKey_184 ^ _zz_CtrlState_nextrndKey_179);
  end

  assign _zz_CtrlState_nextrndKey_185 = (_zz_CtrlState_nextrndKey_168 ^ _zz_CtrlState_nextrndKey_169);
  assign _zz_CtrlState_nextrndKey_188 = _zz_CtrlState_nextrndKey_185[3 : 2];
  assign _zz_CtrlState_nextrndKey_189 = _zz_CtrlState_nextrndKey_185[1 : 0];
  assign _zz_CtrlState_nextrndKey_190 = (_zz_CtrlState_nextrndKey_188 ^ _zz_CtrlState_nextrndKey_189);
  always @(*) begin
    _zz_CtrlState_nextrndKey_191[1] = _zz_CtrlState_nextrndKey_190[1];
    _zz_CtrlState_nextrndKey_191[0] = (_zz_CtrlState_nextrndKey_190[0] ^ _zz_CtrlState_nextrndKey_190[1]);
  end

  assign _zz_CtrlState_nextrndKey_192 = ((_zz_CtrlState_nextrndKey_189[0] && _zz_CtrlState_nextrndKey_188[1]) ^ (_zz_CtrlState_nextrndKey_188[0] && _zz_CtrlState_nextrndKey_189[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_193[1] = ((_zz_CtrlState_nextrndKey_189[0] && _zz_CtrlState_nextrndKey_188[0]) ^ _zz_CtrlState_nextrndKey_192);
    _zz_CtrlState_nextrndKey_193[0] = ((_zz_CtrlState_nextrndKey_189[1] && _zz_CtrlState_nextrndKey_188[1]) ^ _zz_CtrlState_nextrndKey_192);
  end

  assign _zz_CtrlState_nextrndKey_194 = (_zz_CtrlState_nextrndKey_191 ^ _zz_CtrlState_nextrndKey_193);
  always @(*) begin
    _zz_CtrlState_nextrndKey_196[1] = _zz_CtrlState_nextrndKey_194[0];
    _zz_CtrlState_nextrndKey_196[0] = _zz_CtrlState_nextrndKey_194[1];
  end

  assign _zz_CtrlState_nextrndKey_195 = _zz_CtrlState_nextrndKey_196;
  assign _zz_CtrlState_nextrndKey_197 = ((_zz_CtrlState_nextrndKey_195[0] && _zz_CtrlState_nextrndKey_188[1]) ^ (_zz_CtrlState_nextrndKey_188[0] && _zz_CtrlState_nextrndKey_195[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_198[1] = ((_zz_CtrlState_nextrndKey_195[0] && _zz_CtrlState_nextrndKey_188[0]) ^ _zz_CtrlState_nextrndKey_197);
    _zz_CtrlState_nextrndKey_198[0] = ((_zz_CtrlState_nextrndKey_195[1] && _zz_CtrlState_nextrndKey_188[1]) ^ _zz_CtrlState_nextrndKey_197);
  end

  assign _zz_CtrlState_nextrndKey_199 = ((_zz_CtrlState_nextrndKey_195[0] && _zz_CtrlState_nextrndKey_189[1]) ^ (_zz_CtrlState_nextrndKey_189[0] && _zz_CtrlState_nextrndKey_195[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_200[1] = ((_zz_CtrlState_nextrndKey_195[0] && _zz_CtrlState_nextrndKey_189[0]) ^ _zz_CtrlState_nextrndKey_199);
    _zz_CtrlState_nextrndKey_200[0] = ((_zz_CtrlState_nextrndKey_195[1] && _zz_CtrlState_nextrndKey_189[1]) ^ _zz_CtrlState_nextrndKey_199);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_187[3 : 2] = _zz_CtrlState_nextrndKey_200;
    _zz_CtrlState_nextrndKey_187[1 : 0] = _zz_CtrlState_nextrndKey_198;
  end

  assign _zz_CtrlState_nextrndKey_186 = _zz_CtrlState_nextrndKey_187;
  assign _zz_CtrlState_nextrndKey_202 = _zz_CtrlState_nextrndKey_165[3 : 2];
  assign _zz_CtrlState_nextrndKey_203 = _zz_CtrlState_nextrndKey_165[1 : 0];
  assign _zz_CtrlState_nextrndKey_204 = _zz_CtrlState_nextrndKey_186[3 : 2];
  assign _zz_CtrlState_nextrndKey_205 = _zz_CtrlState_nextrndKey_186[1 : 0];
  assign _zz_CtrlState_nextrndKey_206 = (_zz_CtrlState_nextrndKey_202 ^ _zz_CtrlState_nextrndKey_203);
  assign _zz_CtrlState_nextrndKey_207 = (_zz_CtrlState_nextrndKey_204 ^ _zz_CtrlState_nextrndKey_205);
  assign _zz_CtrlState_nextrndKey_209 = ((_zz_CtrlState_nextrndKey_207[0] && _zz_CtrlState_nextrndKey_206[1]) ^ (_zz_CtrlState_nextrndKey_206[0] && _zz_CtrlState_nextrndKey_207[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_210[1] = ((_zz_CtrlState_nextrndKey_207[0] && _zz_CtrlState_nextrndKey_206[0]) ^ _zz_CtrlState_nextrndKey_209);
    _zz_CtrlState_nextrndKey_210[0] = ((_zz_CtrlState_nextrndKey_207[1] && _zz_CtrlState_nextrndKey_206[1]) ^ _zz_CtrlState_nextrndKey_209);
  end

  assign _zz_CtrlState_nextrndKey_208 = _zz_CtrlState_nextrndKey_210;
  always @(*) begin
    _zz_CtrlState_nextrndKey_212[1] = _zz_CtrlState_nextrndKey_208[0];
    _zz_CtrlState_nextrndKey_212[0] = (_zz_CtrlState_nextrndKey_208[0] ^ _zz_CtrlState_nextrndKey_208[1]);
  end

  assign _zz_CtrlState_nextrndKey_211 = _zz_CtrlState_nextrndKey_212;
  assign _zz_CtrlState_nextrndKey_213 = ((_zz_CtrlState_nextrndKey_204[0] && _zz_CtrlState_nextrndKey_202[1]) ^ (_zz_CtrlState_nextrndKey_202[0] && _zz_CtrlState_nextrndKey_204[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_214[1] = ((_zz_CtrlState_nextrndKey_204[0] && _zz_CtrlState_nextrndKey_202[0]) ^ _zz_CtrlState_nextrndKey_213);
    _zz_CtrlState_nextrndKey_214[0] = ((_zz_CtrlState_nextrndKey_204[1] && _zz_CtrlState_nextrndKey_202[1]) ^ _zz_CtrlState_nextrndKey_213);
  end

  assign _zz_CtrlState_nextrndKey_215 = ((_zz_CtrlState_nextrndKey_205[0] && _zz_CtrlState_nextrndKey_203[1]) ^ (_zz_CtrlState_nextrndKey_203[0] && _zz_CtrlState_nextrndKey_205[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_216[1] = ((_zz_CtrlState_nextrndKey_205[0] && _zz_CtrlState_nextrndKey_203[0]) ^ _zz_CtrlState_nextrndKey_215);
    _zz_CtrlState_nextrndKey_216[0] = ((_zz_CtrlState_nextrndKey_205[1] && _zz_CtrlState_nextrndKey_203[1]) ^ _zz_CtrlState_nextrndKey_215);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_201[3 : 2] = (_zz_CtrlState_nextrndKey_214 ^ _zz_CtrlState_nextrndKey_211);
    _zz_CtrlState_nextrndKey_201[1 : 0] = (_zz_CtrlState_nextrndKey_216 ^ _zz_CtrlState_nextrndKey_211);
  end

  assign _zz_CtrlState_nextrndKey_218 = _zz_CtrlState_nextrndKey_166[3 : 2];
  assign _zz_CtrlState_nextrndKey_219 = _zz_CtrlState_nextrndKey_166[1 : 0];
  assign _zz_CtrlState_nextrndKey_220 = _zz_CtrlState_nextrndKey_186[3 : 2];
  assign _zz_CtrlState_nextrndKey_221 = _zz_CtrlState_nextrndKey_186[1 : 0];
  assign _zz_CtrlState_nextrndKey_222 = (_zz_CtrlState_nextrndKey_218 ^ _zz_CtrlState_nextrndKey_219);
  assign _zz_CtrlState_nextrndKey_223 = (_zz_CtrlState_nextrndKey_220 ^ _zz_CtrlState_nextrndKey_221);
  assign _zz_CtrlState_nextrndKey_225 = ((_zz_CtrlState_nextrndKey_223[0] && _zz_CtrlState_nextrndKey_222[1]) ^ (_zz_CtrlState_nextrndKey_222[0] && _zz_CtrlState_nextrndKey_223[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_226[1] = ((_zz_CtrlState_nextrndKey_223[0] && _zz_CtrlState_nextrndKey_222[0]) ^ _zz_CtrlState_nextrndKey_225);
    _zz_CtrlState_nextrndKey_226[0] = ((_zz_CtrlState_nextrndKey_223[1] && _zz_CtrlState_nextrndKey_222[1]) ^ _zz_CtrlState_nextrndKey_225);
  end

  assign _zz_CtrlState_nextrndKey_224 = _zz_CtrlState_nextrndKey_226;
  always @(*) begin
    _zz_CtrlState_nextrndKey_228[1] = _zz_CtrlState_nextrndKey_224[0];
    _zz_CtrlState_nextrndKey_228[0] = (_zz_CtrlState_nextrndKey_224[0] ^ _zz_CtrlState_nextrndKey_224[1]);
  end

  assign _zz_CtrlState_nextrndKey_227 = _zz_CtrlState_nextrndKey_228;
  assign _zz_CtrlState_nextrndKey_229 = ((_zz_CtrlState_nextrndKey_220[0] && _zz_CtrlState_nextrndKey_218[1]) ^ (_zz_CtrlState_nextrndKey_218[0] && _zz_CtrlState_nextrndKey_220[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_230[1] = ((_zz_CtrlState_nextrndKey_220[0] && _zz_CtrlState_nextrndKey_218[0]) ^ _zz_CtrlState_nextrndKey_229);
    _zz_CtrlState_nextrndKey_230[0] = ((_zz_CtrlState_nextrndKey_220[1] && _zz_CtrlState_nextrndKey_218[1]) ^ _zz_CtrlState_nextrndKey_229);
  end

  assign _zz_CtrlState_nextrndKey_231 = ((_zz_CtrlState_nextrndKey_221[0] && _zz_CtrlState_nextrndKey_219[1]) ^ (_zz_CtrlState_nextrndKey_219[0] && _zz_CtrlState_nextrndKey_221[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_232[1] = ((_zz_CtrlState_nextrndKey_221[0] && _zz_CtrlState_nextrndKey_219[0]) ^ _zz_CtrlState_nextrndKey_231);
    _zz_CtrlState_nextrndKey_232[0] = ((_zz_CtrlState_nextrndKey_221[1] && _zz_CtrlState_nextrndKey_219[1]) ^ _zz_CtrlState_nextrndKey_231);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_217[3 : 2] = (_zz_CtrlState_nextrndKey_230 ^ _zz_CtrlState_nextrndKey_227);
    _zz_CtrlState_nextrndKey_217[1 : 0] = (_zz_CtrlState_nextrndKey_232 ^ _zz_CtrlState_nextrndKey_227);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_164[7 : 4] = _zz_CtrlState_nextrndKey_217;
    _zz_CtrlState_nextrndKey_164[3 : 0] = _zz_CtrlState_nextrndKey_201;
  end

  assign _zz_CtrlState_nextrndKey_163 = _zz_CtrlState_nextrndKey_164;
  always @(*) begin
    _zz_CtrlState_nextrndKey_234[7] = (_zz_CtrlState_nextrndKey_163[5] ^ _zz_CtrlState_nextrndKey_163[3]);
    _zz_CtrlState_nextrndKey_234[6] = (_zz_CtrlState_nextrndKey_163[7] ^ _zz_CtrlState_nextrndKey_163[3]);
    _zz_CtrlState_nextrndKey_234[5] = (_zz_CtrlState_nextrndKey_163[6] ^ _zz_CtrlState_nextrndKey_163[0]);
    _zz_CtrlState_nextrndKey_234[4] = ((_zz_CtrlState_nextrndKey_163[7] ^ _zz_CtrlState_nextrndKey_163[5]) ^ _zz_CtrlState_nextrndKey_163[3]);
    _zz_CtrlState_nextrndKey_234[3] = ((((_zz_CtrlState_nextrndKey_163[7] ^ _zz_CtrlState_nextrndKey_163[6]) ^ _zz_CtrlState_nextrndKey_163[5]) ^ _zz_CtrlState_nextrndKey_163[4]) ^ _zz_CtrlState_nextrndKey_163[3]);
    _zz_CtrlState_nextrndKey_234[2] = ((((_zz_CtrlState_nextrndKey_163[6] ^ _zz_CtrlState_nextrndKey_163[5]) ^ _zz_CtrlState_nextrndKey_163[3]) ^ _zz_CtrlState_nextrndKey_163[2]) ^ _zz_CtrlState_nextrndKey_163[0]);
    _zz_CtrlState_nextrndKey_234[1] = ((_zz_CtrlState_nextrndKey_163[5] ^ _zz_CtrlState_nextrndKey_163[4]) ^ _zz_CtrlState_nextrndKey_163[1]);
    _zz_CtrlState_nextrndKey_234[0] = ((_zz_CtrlState_nextrndKey_163[6] ^ _zz_CtrlState_nextrndKey_163[4]) ^ _zz_CtrlState_nextrndKey_163[1]);
  end

  assign _zz_CtrlState_nextrndKey_233 = _zz_CtrlState_nextrndKey_234;
  always @(*) begin
    _zz_CtrlState_nextrndKey_160[7] = _zz_CtrlState_nextrndKey_233[7];
    _zz_CtrlState_nextrndKey_160[6] = (! _zz_CtrlState_nextrndKey_233[6]);
    _zz_CtrlState_nextrndKey_160[5] = (! _zz_CtrlState_nextrndKey_233[5]);
    _zz_CtrlState_nextrndKey_160[4] = _zz_CtrlState_nextrndKey_233[4];
    _zz_CtrlState_nextrndKey_160[3] = _zz_CtrlState_nextrndKey_233[3];
    _zz_CtrlState_nextrndKey_160[2] = _zz_CtrlState_nextrndKey_233[2];
    _zz_CtrlState_nextrndKey_160[1] = (! _zz_CtrlState_nextrndKey_233[1]);
    _zz_CtrlState_nextrndKey_160[0] = (! _zz_CtrlState_nextrndKey_233[0]);
  end

  assign _zz_CtrlState_nextrndKey_235 = _zz_CtrlState_nextrndKey_5[31 : 24];
  always @(*) begin
    _zz_CtrlState_nextrndKey_238[7] = (((((_zz_CtrlState_nextrndKey_235[7] ^ _zz_CtrlState_nextrndKey_235[6]) ^ _zz_CtrlState_nextrndKey_235[5]) ^ _zz_CtrlState_nextrndKey_235[2]) ^ _zz_CtrlState_nextrndKey_235[1]) ^ _zz_CtrlState_nextrndKey_235[0]);
    _zz_CtrlState_nextrndKey_238[6] = (((_zz_CtrlState_nextrndKey_235[6] ^ _zz_CtrlState_nextrndKey_235[5]) ^ _zz_CtrlState_nextrndKey_235[4]) ^ _zz_CtrlState_nextrndKey_235[0]);
    _zz_CtrlState_nextrndKey_238[5] = (((_zz_CtrlState_nextrndKey_235[6] ^ _zz_CtrlState_nextrndKey_235[5]) ^ _zz_CtrlState_nextrndKey_235[1]) ^ _zz_CtrlState_nextrndKey_235[0]);
    _zz_CtrlState_nextrndKey_238[4] = (((_zz_CtrlState_nextrndKey_235[7] ^ _zz_CtrlState_nextrndKey_235[6]) ^ _zz_CtrlState_nextrndKey_235[5]) ^ _zz_CtrlState_nextrndKey_235[0]);
    _zz_CtrlState_nextrndKey_238[3] = ((((_zz_CtrlState_nextrndKey_235[7] ^ _zz_CtrlState_nextrndKey_235[4]) ^ _zz_CtrlState_nextrndKey_235[3]) ^ _zz_CtrlState_nextrndKey_235[1]) ^ _zz_CtrlState_nextrndKey_235[0]);
    _zz_CtrlState_nextrndKey_238[2] = _zz_CtrlState_nextrndKey_235[0];
    _zz_CtrlState_nextrndKey_238[1] = ((_zz_CtrlState_nextrndKey_235[6] ^ _zz_CtrlState_nextrndKey_235[5]) ^ _zz_CtrlState_nextrndKey_235[0]);
    _zz_CtrlState_nextrndKey_238[0] = ((((_zz_CtrlState_nextrndKey_235[6] ^ _zz_CtrlState_nextrndKey_235[3]) ^ _zz_CtrlState_nextrndKey_235[2]) ^ _zz_CtrlState_nextrndKey_235[1]) ^ _zz_CtrlState_nextrndKey_235[0]);
  end

  assign _zz_CtrlState_nextrndKey_237 = _zz_CtrlState_nextrndKey_238;
  assign _zz_CtrlState_nextrndKey_241 = _zz_CtrlState_nextrndKey_237[7 : 4];
  assign _zz_CtrlState_nextrndKey_242 = _zz_CtrlState_nextrndKey_237[3 : 0];
  assign _zz_CtrlState_nextrndKey_243 = (_zz_CtrlState_nextrndKey_241 ^ _zz_CtrlState_nextrndKey_242);
  always @(*) begin
    _zz_CtrlState_nextrndKey_244[3] = (_zz_CtrlState_nextrndKey_243[2] ^ _zz_CtrlState_nextrndKey_243[0]);
    _zz_CtrlState_nextrndKey_244[2] = (_zz_CtrlState_nextrndKey_243[3] ^ _zz_CtrlState_nextrndKey_243[1]);
    _zz_CtrlState_nextrndKey_244[1] = (_zz_CtrlState_nextrndKey_243[1] ^ _zz_CtrlState_nextrndKey_243[0]);
    _zz_CtrlState_nextrndKey_244[0] = _zz_CtrlState_nextrndKey_243[0];
  end

  assign _zz_CtrlState_nextrndKey_246 = _zz_CtrlState_nextrndKey_241[3 : 2];
  assign _zz_CtrlState_nextrndKey_247 = _zz_CtrlState_nextrndKey_241[1 : 0];
  assign _zz_CtrlState_nextrndKey_248 = _zz_CtrlState_nextrndKey_242[3 : 2];
  assign _zz_CtrlState_nextrndKey_249 = _zz_CtrlState_nextrndKey_242[1 : 0];
  assign _zz_CtrlState_nextrndKey_250 = (_zz_CtrlState_nextrndKey_246 ^ _zz_CtrlState_nextrndKey_247);
  assign _zz_CtrlState_nextrndKey_251 = (_zz_CtrlState_nextrndKey_248 ^ _zz_CtrlState_nextrndKey_249);
  assign _zz_CtrlState_nextrndKey_253 = ((_zz_CtrlState_nextrndKey_251[0] && _zz_CtrlState_nextrndKey_250[1]) ^ (_zz_CtrlState_nextrndKey_250[0] && _zz_CtrlState_nextrndKey_251[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_254[1] = ((_zz_CtrlState_nextrndKey_251[0] && _zz_CtrlState_nextrndKey_250[0]) ^ _zz_CtrlState_nextrndKey_253);
    _zz_CtrlState_nextrndKey_254[0] = ((_zz_CtrlState_nextrndKey_251[1] && _zz_CtrlState_nextrndKey_250[1]) ^ _zz_CtrlState_nextrndKey_253);
  end

  assign _zz_CtrlState_nextrndKey_252 = _zz_CtrlState_nextrndKey_254;
  always @(*) begin
    _zz_CtrlState_nextrndKey_256[1] = _zz_CtrlState_nextrndKey_252[0];
    _zz_CtrlState_nextrndKey_256[0] = (_zz_CtrlState_nextrndKey_252[0] ^ _zz_CtrlState_nextrndKey_252[1]);
  end

  assign _zz_CtrlState_nextrndKey_255 = _zz_CtrlState_nextrndKey_256;
  assign _zz_CtrlState_nextrndKey_257 = ((_zz_CtrlState_nextrndKey_248[0] && _zz_CtrlState_nextrndKey_246[1]) ^ (_zz_CtrlState_nextrndKey_246[0] && _zz_CtrlState_nextrndKey_248[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_258[1] = ((_zz_CtrlState_nextrndKey_248[0] && _zz_CtrlState_nextrndKey_246[0]) ^ _zz_CtrlState_nextrndKey_257);
    _zz_CtrlState_nextrndKey_258[0] = ((_zz_CtrlState_nextrndKey_248[1] && _zz_CtrlState_nextrndKey_246[1]) ^ _zz_CtrlState_nextrndKey_257);
  end

  assign _zz_CtrlState_nextrndKey_259 = ((_zz_CtrlState_nextrndKey_249[0] && _zz_CtrlState_nextrndKey_247[1]) ^ (_zz_CtrlState_nextrndKey_247[0] && _zz_CtrlState_nextrndKey_249[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_260[1] = ((_zz_CtrlState_nextrndKey_249[0] && _zz_CtrlState_nextrndKey_247[0]) ^ _zz_CtrlState_nextrndKey_259);
    _zz_CtrlState_nextrndKey_260[0] = ((_zz_CtrlState_nextrndKey_249[1] && _zz_CtrlState_nextrndKey_247[1]) ^ _zz_CtrlState_nextrndKey_259);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_245[3 : 2] = (_zz_CtrlState_nextrndKey_258 ^ _zz_CtrlState_nextrndKey_255);
    _zz_CtrlState_nextrndKey_245[1 : 0] = (_zz_CtrlState_nextrndKey_260 ^ _zz_CtrlState_nextrndKey_255);
  end

  assign _zz_CtrlState_nextrndKey_261 = (_zz_CtrlState_nextrndKey_244 ^ _zz_CtrlState_nextrndKey_245);
  assign _zz_CtrlState_nextrndKey_264 = _zz_CtrlState_nextrndKey_261[3 : 2];
  assign _zz_CtrlState_nextrndKey_265 = _zz_CtrlState_nextrndKey_261[1 : 0];
  assign _zz_CtrlState_nextrndKey_266 = (_zz_CtrlState_nextrndKey_264 ^ _zz_CtrlState_nextrndKey_265);
  always @(*) begin
    _zz_CtrlState_nextrndKey_267[1] = _zz_CtrlState_nextrndKey_266[1];
    _zz_CtrlState_nextrndKey_267[0] = (_zz_CtrlState_nextrndKey_266[0] ^ _zz_CtrlState_nextrndKey_266[1]);
  end

  assign _zz_CtrlState_nextrndKey_268 = ((_zz_CtrlState_nextrndKey_265[0] && _zz_CtrlState_nextrndKey_264[1]) ^ (_zz_CtrlState_nextrndKey_264[0] && _zz_CtrlState_nextrndKey_265[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_269[1] = ((_zz_CtrlState_nextrndKey_265[0] && _zz_CtrlState_nextrndKey_264[0]) ^ _zz_CtrlState_nextrndKey_268);
    _zz_CtrlState_nextrndKey_269[0] = ((_zz_CtrlState_nextrndKey_265[1] && _zz_CtrlState_nextrndKey_264[1]) ^ _zz_CtrlState_nextrndKey_268);
  end

  assign _zz_CtrlState_nextrndKey_270 = (_zz_CtrlState_nextrndKey_267 ^ _zz_CtrlState_nextrndKey_269);
  always @(*) begin
    _zz_CtrlState_nextrndKey_272[1] = _zz_CtrlState_nextrndKey_270[0];
    _zz_CtrlState_nextrndKey_272[0] = _zz_CtrlState_nextrndKey_270[1];
  end

  assign _zz_CtrlState_nextrndKey_271 = _zz_CtrlState_nextrndKey_272;
  assign _zz_CtrlState_nextrndKey_273 = ((_zz_CtrlState_nextrndKey_271[0] && _zz_CtrlState_nextrndKey_264[1]) ^ (_zz_CtrlState_nextrndKey_264[0] && _zz_CtrlState_nextrndKey_271[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_274[1] = ((_zz_CtrlState_nextrndKey_271[0] && _zz_CtrlState_nextrndKey_264[0]) ^ _zz_CtrlState_nextrndKey_273);
    _zz_CtrlState_nextrndKey_274[0] = ((_zz_CtrlState_nextrndKey_271[1] && _zz_CtrlState_nextrndKey_264[1]) ^ _zz_CtrlState_nextrndKey_273);
  end

  assign _zz_CtrlState_nextrndKey_275 = ((_zz_CtrlState_nextrndKey_271[0] && _zz_CtrlState_nextrndKey_265[1]) ^ (_zz_CtrlState_nextrndKey_265[0] && _zz_CtrlState_nextrndKey_271[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_276[1] = ((_zz_CtrlState_nextrndKey_271[0] && _zz_CtrlState_nextrndKey_265[0]) ^ _zz_CtrlState_nextrndKey_275);
    _zz_CtrlState_nextrndKey_276[0] = ((_zz_CtrlState_nextrndKey_271[1] && _zz_CtrlState_nextrndKey_265[1]) ^ _zz_CtrlState_nextrndKey_275);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_263[3 : 2] = _zz_CtrlState_nextrndKey_276;
    _zz_CtrlState_nextrndKey_263[1 : 0] = _zz_CtrlState_nextrndKey_274;
  end

  assign _zz_CtrlState_nextrndKey_262 = _zz_CtrlState_nextrndKey_263;
  assign _zz_CtrlState_nextrndKey_278 = _zz_CtrlState_nextrndKey_241[3 : 2];
  assign _zz_CtrlState_nextrndKey_279 = _zz_CtrlState_nextrndKey_241[1 : 0];
  assign _zz_CtrlState_nextrndKey_280 = _zz_CtrlState_nextrndKey_262[3 : 2];
  assign _zz_CtrlState_nextrndKey_281 = _zz_CtrlState_nextrndKey_262[1 : 0];
  assign _zz_CtrlState_nextrndKey_282 = (_zz_CtrlState_nextrndKey_278 ^ _zz_CtrlState_nextrndKey_279);
  assign _zz_CtrlState_nextrndKey_283 = (_zz_CtrlState_nextrndKey_280 ^ _zz_CtrlState_nextrndKey_281);
  assign _zz_CtrlState_nextrndKey_285 = ((_zz_CtrlState_nextrndKey_283[0] && _zz_CtrlState_nextrndKey_282[1]) ^ (_zz_CtrlState_nextrndKey_282[0] && _zz_CtrlState_nextrndKey_283[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_286[1] = ((_zz_CtrlState_nextrndKey_283[0] && _zz_CtrlState_nextrndKey_282[0]) ^ _zz_CtrlState_nextrndKey_285);
    _zz_CtrlState_nextrndKey_286[0] = ((_zz_CtrlState_nextrndKey_283[1] && _zz_CtrlState_nextrndKey_282[1]) ^ _zz_CtrlState_nextrndKey_285);
  end

  assign _zz_CtrlState_nextrndKey_284 = _zz_CtrlState_nextrndKey_286;
  always @(*) begin
    _zz_CtrlState_nextrndKey_288[1] = _zz_CtrlState_nextrndKey_284[0];
    _zz_CtrlState_nextrndKey_288[0] = (_zz_CtrlState_nextrndKey_284[0] ^ _zz_CtrlState_nextrndKey_284[1]);
  end

  assign _zz_CtrlState_nextrndKey_287 = _zz_CtrlState_nextrndKey_288;
  assign _zz_CtrlState_nextrndKey_289 = ((_zz_CtrlState_nextrndKey_280[0] && _zz_CtrlState_nextrndKey_278[1]) ^ (_zz_CtrlState_nextrndKey_278[0] && _zz_CtrlState_nextrndKey_280[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_290[1] = ((_zz_CtrlState_nextrndKey_280[0] && _zz_CtrlState_nextrndKey_278[0]) ^ _zz_CtrlState_nextrndKey_289);
    _zz_CtrlState_nextrndKey_290[0] = ((_zz_CtrlState_nextrndKey_280[1] && _zz_CtrlState_nextrndKey_278[1]) ^ _zz_CtrlState_nextrndKey_289);
  end

  assign _zz_CtrlState_nextrndKey_291 = ((_zz_CtrlState_nextrndKey_281[0] && _zz_CtrlState_nextrndKey_279[1]) ^ (_zz_CtrlState_nextrndKey_279[0] && _zz_CtrlState_nextrndKey_281[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_292[1] = ((_zz_CtrlState_nextrndKey_281[0] && _zz_CtrlState_nextrndKey_279[0]) ^ _zz_CtrlState_nextrndKey_291);
    _zz_CtrlState_nextrndKey_292[0] = ((_zz_CtrlState_nextrndKey_281[1] && _zz_CtrlState_nextrndKey_279[1]) ^ _zz_CtrlState_nextrndKey_291);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_277[3 : 2] = (_zz_CtrlState_nextrndKey_290 ^ _zz_CtrlState_nextrndKey_287);
    _zz_CtrlState_nextrndKey_277[1 : 0] = (_zz_CtrlState_nextrndKey_292 ^ _zz_CtrlState_nextrndKey_287);
  end

  assign _zz_CtrlState_nextrndKey_294 = _zz_CtrlState_nextrndKey_242[3 : 2];
  assign _zz_CtrlState_nextrndKey_295 = _zz_CtrlState_nextrndKey_242[1 : 0];
  assign _zz_CtrlState_nextrndKey_296 = _zz_CtrlState_nextrndKey_262[3 : 2];
  assign _zz_CtrlState_nextrndKey_297 = _zz_CtrlState_nextrndKey_262[1 : 0];
  assign _zz_CtrlState_nextrndKey_298 = (_zz_CtrlState_nextrndKey_294 ^ _zz_CtrlState_nextrndKey_295);
  assign _zz_CtrlState_nextrndKey_299 = (_zz_CtrlState_nextrndKey_296 ^ _zz_CtrlState_nextrndKey_297);
  assign _zz_CtrlState_nextrndKey_301 = ((_zz_CtrlState_nextrndKey_299[0] && _zz_CtrlState_nextrndKey_298[1]) ^ (_zz_CtrlState_nextrndKey_298[0] && _zz_CtrlState_nextrndKey_299[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_302[1] = ((_zz_CtrlState_nextrndKey_299[0] && _zz_CtrlState_nextrndKey_298[0]) ^ _zz_CtrlState_nextrndKey_301);
    _zz_CtrlState_nextrndKey_302[0] = ((_zz_CtrlState_nextrndKey_299[1] && _zz_CtrlState_nextrndKey_298[1]) ^ _zz_CtrlState_nextrndKey_301);
  end

  assign _zz_CtrlState_nextrndKey_300 = _zz_CtrlState_nextrndKey_302;
  always @(*) begin
    _zz_CtrlState_nextrndKey_304[1] = _zz_CtrlState_nextrndKey_300[0];
    _zz_CtrlState_nextrndKey_304[0] = (_zz_CtrlState_nextrndKey_300[0] ^ _zz_CtrlState_nextrndKey_300[1]);
  end

  assign _zz_CtrlState_nextrndKey_303 = _zz_CtrlState_nextrndKey_304;
  assign _zz_CtrlState_nextrndKey_305 = ((_zz_CtrlState_nextrndKey_296[0] && _zz_CtrlState_nextrndKey_294[1]) ^ (_zz_CtrlState_nextrndKey_294[0] && _zz_CtrlState_nextrndKey_296[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_306[1] = ((_zz_CtrlState_nextrndKey_296[0] && _zz_CtrlState_nextrndKey_294[0]) ^ _zz_CtrlState_nextrndKey_305);
    _zz_CtrlState_nextrndKey_306[0] = ((_zz_CtrlState_nextrndKey_296[1] && _zz_CtrlState_nextrndKey_294[1]) ^ _zz_CtrlState_nextrndKey_305);
  end

  assign _zz_CtrlState_nextrndKey_307 = ((_zz_CtrlState_nextrndKey_297[0] && _zz_CtrlState_nextrndKey_295[1]) ^ (_zz_CtrlState_nextrndKey_295[0] && _zz_CtrlState_nextrndKey_297[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_308[1] = ((_zz_CtrlState_nextrndKey_297[0] && _zz_CtrlState_nextrndKey_295[0]) ^ _zz_CtrlState_nextrndKey_307);
    _zz_CtrlState_nextrndKey_308[0] = ((_zz_CtrlState_nextrndKey_297[1] && _zz_CtrlState_nextrndKey_295[1]) ^ _zz_CtrlState_nextrndKey_307);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_293[3 : 2] = (_zz_CtrlState_nextrndKey_306 ^ _zz_CtrlState_nextrndKey_303);
    _zz_CtrlState_nextrndKey_293[1 : 0] = (_zz_CtrlState_nextrndKey_308 ^ _zz_CtrlState_nextrndKey_303);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_240[7 : 4] = _zz_CtrlState_nextrndKey_293;
    _zz_CtrlState_nextrndKey_240[3 : 0] = _zz_CtrlState_nextrndKey_277;
  end

  assign _zz_CtrlState_nextrndKey_239 = _zz_CtrlState_nextrndKey_240;
  always @(*) begin
    _zz_CtrlState_nextrndKey_310[7] = (_zz_CtrlState_nextrndKey_239[5] ^ _zz_CtrlState_nextrndKey_239[3]);
    _zz_CtrlState_nextrndKey_310[6] = (_zz_CtrlState_nextrndKey_239[7] ^ _zz_CtrlState_nextrndKey_239[3]);
    _zz_CtrlState_nextrndKey_310[5] = (_zz_CtrlState_nextrndKey_239[6] ^ _zz_CtrlState_nextrndKey_239[0]);
    _zz_CtrlState_nextrndKey_310[4] = ((_zz_CtrlState_nextrndKey_239[7] ^ _zz_CtrlState_nextrndKey_239[5]) ^ _zz_CtrlState_nextrndKey_239[3]);
    _zz_CtrlState_nextrndKey_310[3] = ((((_zz_CtrlState_nextrndKey_239[7] ^ _zz_CtrlState_nextrndKey_239[6]) ^ _zz_CtrlState_nextrndKey_239[5]) ^ _zz_CtrlState_nextrndKey_239[4]) ^ _zz_CtrlState_nextrndKey_239[3]);
    _zz_CtrlState_nextrndKey_310[2] = ((((_zz_CtrlState_nextrndKey_239[6] ^ _zz_CtrlState_nextrndKey_239[5]) ^ _zz_CtrlState_nextrndKey_239[3]) ^ _zz_CtrlState_nextrndKey_239[2]) ^ _zz_CtrlState_nextrndKey_239[0]);
    _zz_CtrlState_nextrndKey_310[1] = ((_zz_CtrlState_nextrndKey_239[5] ^ _zz_CtrlState_nextrndKey_239[4]) ^ _zz_CtrlState_nextrndKey_239[1]);
    _zz_CtrlState_nextrndKey_310[0] = ((_zz_CtrlState_nextrndKey_239[6] ^ _zz_CtrlState_nextrndKey_239[4]) ^ _zz_CtrlState_nextrndKey_239[1]);
  end

  assign _zz_CtrlState_nextrndKey_309 = _zz_CtrlState_nextrndKey_310;
  always @(*) begin
    _zz_CtrlState_nextrndKey_236[7] = _zz_CtrlState_nextrndKey_309[7];
    _zz_CtrlState_nextrndKey_236[6] = (! _zz_CtrlState_nextrndKey_309[6]);
    _zz_CtrlState_nextrndKey_236[5] = (! _zz_CtrlState_nextrndKey_309[5]);
    _zz_CtrlState_nextrndKey_236[4] = _zz_CtrlState_nextrndKey_309[4];
    _zz_CtrlState_nextrndKey_236[3] = _zz_CtrlState_nextrndKey_309[3];
    _zz_CtrlState_nextrndKey_236[2] = _zz_CtrlState_nextrndKey_309[2];
    _zz_CtrlState_nextrndKey_236[1] = (! _zz_CtrlState_nextrndKey_309[1]);
    _zz_CtrlState_nextrndKey_236[0] = (! _zz_CtrlState_nextrndKey_309[0]);
  end

  assign _zz_CtrlState_nextrndKey_1 = (_zz_CtrlState_nextrndKey[31 : 0] ^ {(_zz_CtrlState_nextrndKey_6[31 : 24] ^ 8'h01),{_zz_CtrlState_nextrndKey_6[23 : 16],{_zz_CtrlState_nextrndKey_6[15 : 8],_zz_CtrlState_nextrndKey_6[7 : 0]}}});
  assign _zz_CtrlState_nextrndKey_2 = (_zz_CtrlState_nextrndKey[63 : 32] ^ _zz_CtrlState_nextrndKey_1);
  assign _zz_CtrlState_nextrndKey_3 = (_zz_CtrlState_nextrndKey[95 : 64] ^ _zz_CtrlState_nextrndKey_2);
  assign _zz_CtrlState_nextrndKey_311 = {CtrlState_nextrndKey[31 : 0],{CtrlState_nextrndKey[63 : 32],{CtrlState_nextrndKey[95 : 64],CtrlState_nextrndKey[127 : 96]}}};
  assign _zz_CtrlState_nextrndKey_312 = (CtrlState_rndCnt + 4'b0001);
  assign _zz_CtrlState_nextrndKey_316 = _zz_CtrlState_nextrndKey_311[127 : 96];
  assign _zz_CtrlState_nextrndKey_317 = {_zz_CtrlState_nextrndKey_316[23 : 0],_zz_CtrlState_nextrndKey_316[31 : 24]};
  assign _zz_CtrlState_nextrndKey_319 = _zz_CtrlState_nextrndKey_317[7 : 0];
  always @(*) begin
    _zz_CtrlState_nextrndKey_322[7] = (((((_zz_CtrlState_nextrndKey_319[7] ^ _zz_CtrlState_nextrndKey_319[6]) ^ _zz_CtrlState_nextrndKey_319[5]) ^ _zz_CtrlState_nextrndKey_319[2]) ^ _zz_CtrlState_nextrndKey_319[1]) ^ _zz_CtrlState_nextrndKey_319[0]);
    _zz_CtrlState_nextrndKey_322[6] = (((_zz_CtrlState_nextrndKey_319[6] ^ _zz_CtrlState_nextrndKey_319[5]) ^ _zz_CtrlState_nextrndKey_319[4]) ^ _zz_CtrlState_nextrndKey_319[0]);
    _zz_CtrlState_nextrndKey_322[5] = (((_zz_CtrlState_nextrndKey_319[6] ^ _zz_CtrlState_nextrndKey_319[5]) ^ _zz_CtrlState_nextrndKey_319[1]) ^ _zz_CtrlState_nextrndKey_319[0]);
    _zz_CtrlState_nextrndKey_322[4] = (((_zz_CtrlState_nextrndKey_319[7] ^ _zz_CtrlState_nextrndKey_319[6]) ^ _zz_CtrlState_nextrndKey_319[5]) ^ _zz_CtrlState_nextrndKey_319[0]);
    _zz_CtrlState_nextrndKey_322[3] = ((((_zz_CtrlState_nextrndKey_319[7] ^ _zz_CtrlState_nextrndKey_319[4]) ^ _zz_CtrlState_nextrndKey_319[3]) ^ _zz_CtrlState_nextrndKey_319[1]) ^ _zz_CtrlState_nextrndKey_319[0]);
    _zz_CtrlState_nextrndKey_322[2] = _zz_CtrlState_nextrndKey_319[0];
    _zz_CtrlState_nextrndKey_322[1] = ((_zz_CtrlState_nextrndKey_319[6] ^ _zz_CtrlState_nextrndKey_319[5]) ^ _zz_CtrlState_nextrndKey_319[0]);
    _zz_CtrlState_nextrndKey_322[0] = ((((_zz_CtrlState_nextrndKey_319[6] ^ _zz_CtrlState_nextrndKey_319[3]) ^ _zz_CtrlState_nextrndKey_319[2]) ^ _zz_CtrlState_nextrndKey_319[1]) ^ _zz_CtrlState_nextrndKey_319[0]);
  end

  assign _zz_CtrlState_nextrndKey_321 = _zz_CtrlState_nextrndKey_322;
  assign _zz_CtrlState_nextrndKey_325 = _zz_CtrlState_nextrndKey_321[7 : 4];
  assign _zz_CtrlState_nextrndKey_326 = _zz_CtrlState_nextrndKey_321[3 : 0];
  assign _zz_CtrlState_nextrndKey_327 = (_zz_CtrlState_nextrndKey_325 ^ _zz_CtrlState_nextrndKey_326);
  always @(*) begin
    _zz_CtrlState_nextrndKey_328[3] = (_zz_CtrlState_nextrndKey_327[2] ^ _zz_CtrlState_nextrndKey_327[0]);
    _zz_CtrlState_nextrndKey_328[2] = (_zz_CtrlState_nextrndKey_327[3] ^ _zz_CtrlState_nextrndKey_327[1]);
    _zz_CtrlState_nextrndKey_328[1] = (_zz_CtrlState_nextrndKey_327[1] ^ _zz_CtrlState_nextrndKey_327[0]);
    _zz_CtrlState_nextrndKey_328[0] = _zz_CtrlState_nextrndKey_327[0];
  end

  assign _zz_CtrlState_nextrndKey_330 = _zz_CtrlState_nextrndKey_325[3 : 2];
  assign _zz_CtrlState_nextrndKey_331 = _zz_CtrlState_nextrndKey_325[1 : 0];
  assign _zz_CtrlState_nextrndKey_332 = _zz_CtrlState_nextrndKey_326[3 : 2];
  assign _zz_CtrlState_nextrndKey_333 = _zz_CtrlState_nextrndKey_326[1 : 0];
  assign _zz_CtrlState_nextrndKey_334 = (_zz_CtrlState_nextrndKey_330 ^ _zz_CtrlState_nextrndKey_331);
  assign _zz_CtrlState_nextrndKey_335 = (_zz_CtrlState_nextrndKey_332 ^ _zz_CtrlState_nextrndKey_333);
  assign _zz_CtrlState_nextrndKey_337 = ((_zz_CtrlState_nextrndKey_335[0] && _zz_CtrlState_nextrndKey_334[1]) ^ (_zz_CtrlState_nextrndKey_334[0] && _zz_CtrlState_nextrndKey_335[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_338[1] = ((_zz_CtrlState_nextrndKey_335[0] && _zz_CtrlState_nextrndKey_334[0]) ^ _zz_CtrlState_nextrndKey_337);
    _zz_CtrlState_nextrndKey_338[0] = ((_zz_CtrlState_nextrndKey_335[1] && _zz_CtrlState_nextrndKey_334[1]) ^ _zz_CtrlState_nextrndKey_337);
  end

  assign _zz_CtrlState_nextrndKey_336 = _zz_CtrlState_nextrndKey_338;
  always @(*) begin
    _zz_CtrlState_nextrndKey_340[1] = _zz_CtrlState_nextrndKey_336[0];
    _zz_CtrlState_nextrndKey_340[0] = (_zz_CtrlState_nextrndKey_336[0] ^ _zz_CtrlState_nextrndKey_336[1]);
  end

  assign _zz_CtrlState_nextrndKey_339 = _zz_CtrlState_nextrndKey_340;
  assign _zz_CtrlState_nextrndKey_341 = ((_zz_CtrlState_nextrndKey_332[0] && _zz_CtrlState_nextrndKey_330[1]) ^ (_zz_CtrlState_nextrndKey_330[0] && _zz_CtrlState_nextrndKey_332[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_342[1] = ((_zz_CtrlState_nextrndKey_332[0] && _zz_CtrlState_nextrndKey_330[0]) ^ _zz_CtrlState_nextrndKey_341);
    _zz_CtrlState_nextrndKey_342[0] = ((_zz_CtrlState_nextrndKey_332[1] && _zz_CtrlState_nextrndKey_330[1]) ^ _zz_CtrlState_nextrndKey_341);
  end

  assign _zz_CtrlState_nextrndKey_343 = ((_zz_CtrlState_nextrndKey_333[0] && _zz_CtrlState_nextrndKey_331[1]) ^ (_zz_CtrlState_nextrndKey_331[0] && _zz_CtrlState_nextrndKey_333[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_344[1] = ((_zz_CtrlState_nextrndKey_333[0] && _zz_CtrlState_nextrndKey_331[0]) ^ _zz_CtrlState_nextrndKey_343);
    _zz_CtrlState_nextrndKey_344[0] = ((_zz_CtrlState_nextrndKey_333[1] && _zz_CtrlState_nextrndKey_331[1]) ^ _zz_CtrlState_nextrndKey_343);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_329[3 : 2] = (_zz_CtrlState_nextrndKey_342 ^ _zz_CtrlState_nextrndKey_339);
    _zz_CtrlState_nextrndKey_329[1 : 0] = (_zz_CtrlState_nextrndKey_344 ^ _zz_CtrlState_nextrndKey_339);
  end

  assign _zz_CtrlState_nextrndKey_345 = (_zz_CtrlState_nextrndKey_328 ^ _zz_CtrlState_nextrndKey_329);
  assign _zz_CtrlState_nextrndKey_348 = _zz_CtrlState_nextrndKey_345[3 : 2];
  assign _zz_CtrlState_nextrndKey_349 = _zz_CtrlState_nextrndKey_345[1 : 0];
  assign _zz_CtrlState_nextrndKey_350 = (_zz_CtrlState_nextrndKey_348 ^ _zz_CtrlState_nextrndKey_349);
  always @(*) begin
    _zz_CtrlState_nextrndKey_351[1] = _zz_CtrlState_nextrndKey_350[1];
    _zz_CtrlState_nextrndKey_351[0] = (_zz_CtrlState_nextrndKey_350[0] ^ _zz_CtrlState_nextrndKey_350[1]);
  end

  assign _zz_CtrlState_nextrndKey_352 = ((_zz_CtrlState_nextrndKey_349[0] && _zz_CtrlState_nextrndKey_348[1]) ^ (_zz_CtrlState_nextrndKey_348[0] && _zz_CtrlState_nextrndKey_349[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_353[1] = ((_zz_CtrlState_nextrndKey_349[0] && _zz_CtrlState_nextrndKey_348[0]) ^ _zz_CtrlState_nextrndKey_352);
    _zz_CtrlState_nextrndKey_353[0] = ((_zz_CtrlState_nextrndKey_349[1] && _zz_CtrlState_nextrndKey_348[1]) ^ _zz_CtrlState_nextrndKey_352);
  end

  assign _zz_CtrlState_nextrndKey_354 = (_zz_CtrlState_nextrndKey_351 ^ _zz_CtrlState_nextrndKey_353);
  always @(*) begin
    _zz_CtrlState_nextrndKey_356[1] = _zz_CtrlState_nextrndKey_354[0];
    _zz_CtrlState_nextrndKey_356[0] = _zz_CtrlState_nextrndKey_354[1];
  end

  assign _zz_CtrlState_nextrndKey_355 = _zz_CtrlState_nextrndKey_356;
  assign _zz_CtrlState_nextrndKey_357 = ((_zz_CtrlState_nextrndKey_355[0] && _zz_CtrlState_nextrndKey_348[1]) ^ (_zz_CtrlState_nextrndKey_348[0] && _zz_CtrlState_nextrndKey_355[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_358[1] = ((_zz_CtrlState_nextrndKey_355[0] && _zz_CtrlState_nextrndKey_348[0]) ^ _zz_CtrlState_nextrndKey_357);
    _zz_CtrlState_nextrndKey_358[0] = ((_zz_CtrlState_nextrndKey_355[1] && _zz_CtrlState_nextrndKey_348[1]) ^ _zz_CtrlState_nextrndKey_357);
  end

  assign _zz_CtrlState_nextrndKey_359 = ((_zz_CtrlState_nextrndKey_355[0] && _zz_CtrlState_nextrndKey_349[1]) ^ (_zz_CtrlState_nextrndKey_349[0] && _zz_CtrlState_nextrndKey_355[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_360[1] = ((_zz_CtrlState_nextrndKey_355[0] && _zz_CtrlState_nextrndKey_349[0]) ^ _zz_CtrlState_nextrndKey_359);
    _zz_CtrlState_nextrndKey_360[0] = ((_zz_CtrlState_nextrndKey_355[1] && _zz_CtrlState_nextrndKey_349[1]) ^ _zz_CtrlState_nextrndKey_359);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_347[3 : 2] = _zz_CtrlState_nextrndKey_360;
    _zz_CtrlState_nextrndKey_347[1 : 0] = _zz_CtrlState_nextrndKey_358;
  end

  assign _zz_CtrlState_nextrndKey_346 = _zz_CtrlState_nextrndKey_347;
  assign _zz_CtrlState_nextrndKey_362 = _zz_CtrlState_nextrndKey_325[3 : 2];
  assign _zz_CtrlState_nextrndKey_363 = _zz_CtrlState_nextrndKey_325[1 : 0];
  assign _zz_CtrlState_nextrndKey_364 = _zz_CtrlState_nextrndKey_346[3 : 2];
  assign _zz_CtrlState_nextrndKey_365 = _zz_CtrlState_nextrndKey_346[1 : 0];
  assign _zz_CtrlState_nextrndKey_366 = (_zz_CtrlState_nextrndKey_362 ^ _zz_CtrlState_nextrndKey_363);
  assign _zz_CtrlState_nextrndKey_367 = (_zz_CtrlState_nextrndKey_364 ^ _zz_CtrlState_nextrndKey_365);
  assign _zz_CtrlState_nextrndKey_369 = ((_zz_CtrlState_nextrndKey_367[0] && _zz_CtrlState_nextrndKey_366[1]) ^ (_zz_CtrlState_nextrndKey_366[0] && _zz_CtrlState_nextrndKey_367[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_370[1] = ((_zz_CtrlState_nextrndKey_367[0] && _zz_CtrlState_nextrndKey_366[0]) ^ _zz_CtrlState_nextrndKey_369);
    _zz_CtrlState_nextrndKey_370[0] = ((_zz_CtrlState_nextrndKey_367[1] && _zz_CtrlState_nextrndKey_366[1]) ^ _zz_CtrlState_nextrndKey_369);
  end

  assign _zz_CtrlState_nextrndKey_368 = _zz_CtrlState_nextrndKey_370;
  always @(*) begin
    _zz_CtrlState_nextrndKey_372[1] = _zz_CtrlState_nextrndKey_368[0];
    _zz_CtrlState_nextrndKey_372[0] = (_zz_CtrlState_nextrndKey_368[0] ^ _zz_CtrlState_nextrndKey_368[1]);
  end

  assign _zz_CtrlState_nextrndKey_371 = _zz_CtrlState_nextrndKey_372;
  assign _zz_CtrlState_nextrndKey_373 = ((_zz_CtrlState_nextrndKey_364[0] && _zz_CtrlState_nextrndKey_362[1]) ^ (_zz_CtrlState_nextrndKey_362[0] && _zz_CtrlState_nextrndKey_364[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_374[1] = ((_zz_CtrlState_nextrndKey_364[0] && _zz_CtrlState_nextrndKey_362[0]) ^ _zz_CtrlState_nextrndKey_373);
    _zz_CtrlState_nextrndKey_374[0] = ((_zz_CtrlState_nextrndKey_364[1] && _zz_CtrlState_nextrndKey_362[1]) ^ _zz_CtrlState_nextrndKey_373);
  end

  assign _zz_CtrlState_nextrndKey_375 = ((_zz_CtrlState_nextrndKey_365[0] && _zz_CtrlState_nextrndKey_363[1]) ^ (_zz_CtrlState_nextrndKey_363[0] && _zz_CtrlState_nextrndKey_365[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_376[1] = ((_zz_CtrlState_nextrndKey_365[0] && _zz_CtrlState_nextrndKey_363[0]) ^ _zz_CtrlState_nextrndKey_375);
    _zz_CtrlState_nextrndKey_376[0] = ((_zz_CtrlState_nextrndKey_365[1] && _zz_CtrlState_nextrndKey_363[1]) ^ _zz_CtrlState_nextrndKey_375);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_361[3 : 2] = (_zz_CtrlState_nextrndKey_374 ^ _zz_CtrlState_nextrndKey_371);
    _zz_CtrlState_nextrndKey_361[1 : 0] = (_zz_CtrlState_nextrndKey_376 ^ _zz_CtrlState_nextrndKey_371);
  end

  assign _zz_CtrlState_nextrndKey_378 = _zz_CtrlState_nextrndKey_326[3 : 2];
  assign _zz_CtrlState_nextrndKey_379 = _zz_CtrlState_nextrndKey_326[1 : 0];
  assign _zz_CtrlState_nextrndKey_380 = _zz_CtrlState_nextrndKey_346[3 : 2];
  assign _zz_CtrlState_nextrndKey_381 = _zz_CtrlState_nextrndKey_346[1 : 0];
  assign _zz_CtrlState_nextrndKey_382 = (_zz_CtrlState_nextrndKey_378 ^ _zz_CtrlState_nextrndKey_379);
  assign _zz_CtrlState_nextrndKey_383 = (_zz_CtrlState_nextrndKey_380 ^ _zz_CtrlState_nextrndKey_381);
  assign _zz_CtrlState_nextrndKey_385 = ((_zz_CtrlState_nextrndKey_383[0] && _zz_CtrlState_nextrndKey_382[1]) ^ (_zz_CtrlState_nextrndKey_382[0] && _zz_CtrlState_nextrndKey_383[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_386[1] = ((_zz_CtrlState_nextrndKey_383[0] && _zz_CtrlState_nextrndKey_382[0]) ^ _zz_CtrlState_nextrndKey_385);
    _zz_CtrlState_nextrndKey_386[0] = ((_zz_CtrlState_nextrndKey_383[1] && _zz_CtrlState_nextrndKey_382[1]) ^ _zz_CtrlState_nextrndKey_385);
  end

  assign _zz_CtrlState_nextrndKey_384 = _zz_CtrlState_nextrndKey_386;
  always @(*) begin
    _zz_CtrlState_nextrndKey_388[1] = _zz_CtrlState_nextrndKey_384[0];
    _zz_CtrlState_nextrndKey_388[0] = (_zz_CtrlState_nextrndKey_384[0] ^ _zz_CtrlState_nextrndKey_384[1]);
  end

  assign _zz_CtrlState_nextrndKey_387 = _zz_CtrlState_nextrndKey_388;
  assign _zz_CtrlState_nextrndKey_389 = ((_zz_CtrlState_nextrndKey_380[0] && _zz_CtrlState_nextrndKey_378[1]) ^ (_zz_CtrlState_nextrndKey_378[0] && _zz_CtrlState_nextrndKey_380[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_390[1] = ((_zz_CtrlState_nextrndKey_380[0] && _zz_CtrlState_nextrndKey_378[0]) ^ _zz_CtrlState_nextrndKey_389);
    _zz_CtrlState_nextrndKey_390[0] = ((_zz_CtrlState_nextrndKey_380[1] && _zz_CtrlState_nextrndKey_378[1]) ^ _zz_CtrlState_nextrndKey_389);
  end

  assign _zz_CtrlState_nextrndKey_391 = ((_zz_CtrlState_nextrndKey_381[0] && _zz_CtrlState_nextrndKey_379[1]) ^ (_zz_CtrlState_nextrndKey_379[0] && _zz_CtrlState_nextrndKey_381[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_392[1] = ((_zz_CtrlState_nextrndKey_381[0] && _zz_CtrlState_nextrndKey_379[0]) ^ _zz_CtrlState_nextrndKey_391);
    _zz_CtrlState_nextrndKey_392[0] = ((_zz_CtrlState_nextrndKey_381[1] && _zz_CtrlState_nextrndKey_379[1]) ^ _zz_CtrlState_nextrndKey_391);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_377[3 : 2] = (_zz_CtrlState_nextrndKey_390 ^ _zz_CtrlState_nextrndKey_387);
    _zz_CtrlState_nextrndKey_377[1 : 0] = (_zz_CtrlState_nextrndKey_392 ^ _zz_CtrlState_nextrndKey_387);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_324[7 : 4] = _zz_CtrlState_nextrndKey_377;
    _zz_CtrlState_nextrndKey_324[3 : 0] = _zz_CtrlState_nextrndKey_361;
  end

  assign _zz_CtrlState_nextrndKey_323 = _zz_CtrlState_nextrndKey_324;
  always @(*) begin
    _zz_CtrlState_nextrndKey_394[7] = (_zz_CtrlState_nextrndKey_323[5] ^ _zz_CtrlState_nextrndKey_323[3]);
    _zz_CtrlState_nextrndKey_394[6] = (_zz_CtrlState_nextrndKey_323[7] ^ _zz_CtrlState_nextrndKey_323[3]);
    _zz_CtrlState_nextrndKey_394[5] = (_zz_CtrlState_nextrndKey_323[6] ^ _zz_CtrlState_nextrndKey_323[0]);
    _zz_CtrlState_nextrndKey_394[4] = ((_zz_CtrlState_nextrndKey_323[7] ^ _zz_CtrlState_nextrndKey_323[5]) ^ _zz_CtrlState_nextrndKey_323[3]);
    _zz_CtrlState_nextrndKey_394[3] = ((((_zz_CtrlState_nextrndKey_323[7] ^ _zz_CtrlState_nextrndKey_323[6]) ^ _zz_CtrlState_nextrndKey_323[5]) ^ _zz_CtrlState_nextrndKey_323[4]) ^ _zz_CtrlState_nextrndKey_323[3]);
    _zz_CtrlState_nextrndKey_394[2] = ((((_zz_CtrlState_nextrndKey_323[6] ^ _zz_CtrlState_nextrndKey_323[5]) ^ _zz_CtrlState_nextrndKey_323[3]) ^ _zz_CtrlState_nextrndKey_323[2]) ^ _zz_CtrlState_nextrndKey_323[0]);
    _zz_CtrlState_nextrndKey_394[1] = ((_zz_CtrlState_nextrndKey_323[5] ^ _zz_CtrlState_nextrndKey_323[4]) ^ _zz_CtrlState_nextrndKey_323[1]);
    _zz_CtrlState_nextrndKey_394[0] = ((_zz_CtrlState_nextrndKey_323[6] ^ _zz_CtrlState_nextrndKey_323[4]) ^ _zz_CtrlState_nextrndKey_323[1]);
  end

  assign _zz_CtrlState_nextrndKey_393 = _zz_CtrlState_nextrndKey_394;
  always @(*) begin
    _zz_CtrlState_nextrndKey_320[7] = _zz_CtrlState_nextrndKey_393[7];
    _zz_CtrlState_nextrndKey_320[6] = (! _zz_CtrlState_nextrndKey_393[6]);
    _zz_CtrlState_nextrndKey_320[5] = (! _zz_CtrlState_nextrndKey_393[5]);
    _zz_CtrlState_nextrndKey_320[4] = _zz_CtrlState_nextrndKey_393[4];
    _zz_CtrlState_nextrndKey_320[3] = _zz_CtrlState_nextrndKey_393[3];
    _zz_CtrlState_nextrndKey_320[2] = _zz_CtrlState_nextrndKey_393[2];
    _zz_CtrlState_nextrndKey_320[1] = (! _zz_CtrlState_nextrndKey_393[1]);
    _zz_CtrlState_nextrndKey_320[0] = (! _zz_CtrlState_nextrndKey_393[0]);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_318[7 : 0] = _zz_CtrlState_nextrndKey_320;
    _zz_CtrlState_nextrndKey_318[15 : 8] = _zz_CtrlState_nextrndKey_396;
    _zz_CtrlState_nextrndKey_318[23 : 16] = _zz_CtrlState_nextrndKey_472;
    _zz_CtrlState_nextrndKey_318[31 : 24] = _zz_CtrlState_nextrndKey_548;
  end

  assign _zz_CtrlState_nextrndKey_395 = _zz_CtrlState_nextrndKey_317[15 : 8];
  always @(*) begin
    _zz_CtrlState_nextrndKey_398[7] = (((((_zz_CtrlState_nextrndKey_395[7] ^ _zz_CtrlState_nextrndKey_395[6]) ^ _zz_CtrlState_nextrndKey_395[5]) ^ _zz_CtrlState_nextrndKey_395[2]) ^ _zz_CtrlState_nextrndKey_395[1]) ^ _zz_CtrlState_nextrndKey_395[0]);
    _zz_CtrlState_nextrndKey_398[6] = (((_zz_CtrlState_nextrndKey_395[6] ^ _zz_CtrlState_nextrndKey_395[5]) ^ _zz_CtrlState_nextrndKey_395[4]) ^ _zz_CtrlState_nextrndKey_395[0]);
    _zz_CtrlState_nextrndKey_398[5] = (((_zz_CtrlState_nextrndKey_395[6] ^ _zz_CtrlState_nextrndKey_395[5]) ^ _zz_CtrlState_nextrndKey_395[1]) ^ _zz_CtrlState_nextrndKey_395[0]);
    _zz_CtrlState_nextrndKey_398[4] = (((_zz_CtrlState_nextrndKey_395[7] ^ _zz_CtrlState_nextrndKey_395[6]) ^ _zz_CtrlState_nextrndKey_395[5]) ^ _zz_CtrlState_nextrndKey_395[0]);
    _zz_CtrlState_nextrndKey_398[3] = ((((_zz_CtrlState_nextrndKey_395[7] ^ _zz_CtrlState_nextrndKey_395[4]) ^ _zz_CtrlState_nextrndKey_395[3]) ^ _zz_CtrlState_nextrndKey_395[1]) ^ _zz_CtrlState_nextrndKey_395[0]);
    _zz_CtrlState_nextrndKey_398[2] = _zz_CtrlState_nextrndKey_395[0];
    _zz_CtrlState_nextrndKey_398[1] = ((_zz_CtrlState_nextrndKey_395[6] ^ _zz_CtrlState_nextrndKey_395[5]) ^ _zz_CtrlState_nextrndKey_395[0]);
    _zz_CtrlState_nextrndKey_398[0] = ((((_zz_CtrlState_nextrndKey_395[6] ^ _zz_CtrlState_nextrndKey_395[3]) ^ _zz_CtrlState_nextrndKey_395[2]) ^ _zz_CtrlState_nextrndKey_395[1]) ^ _zz_CtrlState_nextrndKey_395[0]);
  end

  assign _zz_CtrlState_nextrndKey_397 = _zz_CtrlState_nextrndKey_398;
  assign _zz_CtrlState_nextrndKey_401 = _zz_CtrlState_nextrndKey_397[7 : 4];
  assign _zz_CtrlState_nextrndKey_402 = _zz_CtrlState_nextrndKey_397[3 : 0];
  assign _zz_CtrlState_nextrndKey_403 = (_zz_CtrlState_nextrndKey_401 ^ _zz_CtrlState_nextrndKey_402);
  always @(*) begin
    _zz_CtrlState_nextrndKey_404[3] = (_zz_CtrlState_nextrndKey_403[2] ^ _zz_CtrlState_nextrndKey_403[0]);
    _zz_CtrlState_nextrndKey_404[2] = (_zz_CtrlState_nextrndKey_403[3] ^ _zz_CtrlState_nextrndKey_403[1]);
    _zz_CtrlState_nextrndKey_404[1] = (_zz_CtrlState_nextrndKey_403[1] ^ _zz_CtrlState_nextrndKey_403[0]);
    _zz_CtrlState_nextrndKey_404[0] = _zz_CtrlState_nextrndKey_403[0];
  end

  assign _zz_CtrlState_nextrndKey_406 = _zz_CtrlState_nextrndKey_401[3 : 2];
  assign _zz_CtrlState_nextrndKey_407 = _zz_CtrlState_nextrndKey_401[1 : 0];
  assign _zz_CtrlState_nextrndKey_408 = _zz_CtrlState_nextrndKey_402[3 : 2];
  assign _zz_CtrlState_nextrndKey_409 = _zz_CtrlState_nextrndKey_402[1 : 0];
  assign _zz_CtrlState_nextrndKey_410 = (_zz_CtrlState_nextrndKey_406 ^ _zz_CtrlState_nextrndKey_407);
  assign _zz_CtrlState_nextrndKey_411 = (_zz_CtrlState_nextrndKey_408 ^ _zz_CtrlState_nextrndKey_409);
  assign _zz_CtrlState_nextrndKey_413 = ((_zz_CtrlState_nextrndKey_411[0] && _zz_CtrlState_nextrndKey_410[1]) ^ (_zz_CtrlState_nextrndKey_410[0] && _zz_CtrlState_nextrndKey_411[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_414[1] = ((_zz_CtrlState_nextrndKey_411[0] && _zz_CtrlState_nextrndKey_410[0]) ^ _zz_CtrlState_nextrndKey_413);
    _zz_CtrlState_nextrndKey_414[0] = ((_zz_CtrlState_nextrndKey_411[1] && _zz_CtrlState_nextrndKey_410[1]) ^ _zz_CtrlState_nextrndKey_413);
  end

  assign _zz_CtrlState_nextrndKey_412 = _zz_CtrlState_nextrndKey_414;
  always @(*) begin
    _zz_CtrlState_nextrndKey_416[1] = _zz_CtrlState_nextrndKey_412[0];
    _zz_CtrlState_nextrndKey_416[0] = (_zz_CtrlState_nextrndKey_412[0] ^ _zz_CtrlState_nextrndKey_412[1]);
  end

  assign _zz_CtrlState_nextrndKey_415 = _zz_CtrlState_nextrndKey_416;
  assign _zz_CtrlState_nextrndKey_417 = ((_zz_CtrlState_nextrndKey_408[0] && _zz_CtrlState_nextrndKey_406[1]) ^ (_zz_CtrlState_nextrndKey_406[0] && _zz_CtrlState_nextrndKey_408[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_418[1] = ((_zz_CtrlState_nextrndKey_408[0] && _zz_CtrlState_nextrndKey_406[0]) ^ _zz_CtrlState_nextrndKey_417);
    _zz_CtrlState_nextrndKey_418[0] = ((_zz_CtrlState_nextrndKey_408[1] && _zz_CtrlState_nextrndKey_406[1]) ^ _zz_CtrlState_nextrndKey_417);
  end

  assign _zz_CtrlState_nextrndKey_419 = ((_zz_CtrlState_nextrndKey_409[0] && _zz_CtrlState_nextrndKey_407[1]) ^ (_zz_CtrlState_nextrndKey_407[0] && _zz_CtrlState_nextrndKey_409[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_420[1] = ((_zz_CtrlState_nextrndKey_409[0] && _zz_CtrlState_nextrndKey_407[0]) ^ _zz_CtrlState_nextrndKey_419);
    _zz_CtrlState_nextrndKey_420[0] = ((_zz_CtrlState_nextrndKey_409[1] && _zz_CtrlState_nextrndKey_407[1]) ^ _zz_CtrlState_nextrndKey_419);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_405[3 : 2] = (_zz_CtrlState_nextrndKey_418 ^ _zz_CtrlState_nextrndKey_415);
    _zz_CtrlState_nextrndKey_405[1 : 0] = (_zz_CtrlState_nextrndKey_420 ^ _zz_CtrlState_nextrndKey_415);
  end

  assign _zz_CtrlState_nextrndKey_421 = (_zz_CtrlState_nextrndKey_404 ^ _zz_CtrlState_nextrndKey_405);
  assign _zz_CtrlState_nextrndKey_424 = _zz_CtrlState_nextrndKey_421[3 : 2];
  assign _zz_CtrlState_nextrndKey_425 = _zz_CtrlState_nextrndKey_421[1 : 0];
  assign _zz_CtrlState_nextrndKey_426 = (_zz_CtrlState_nextrndKey_424 ^ _zz_CtrlState_nextrndKey_425);
  always @(*) begin
    _zz_CtrlState_nextrndKey_427[1] = _zz_CtrlState_nextrndKey_426[1];
    _zz_CtrlState_nextrndKey_427[0] = (_zz_CtrlState_nextrndKey_426[0] ^ _zz_CtrlState_nextrndKey_426[1]);
  end

  assign _zz_CtrlState_nextrndKey_428 = ((_zz_CtrlState_nextrndKey_425[0] && _zz_CtrlState_nextrndKey_424[1]) ^ (_zz_CtrlState_nextrndKey_424[0] && _zz_CtrlState_nextrndKey_425[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_429[1] = ((_zz_CtrlState_nextrndKey_425[0] && _zz_CtrlState_nextrndKey_424[0]) ^ _zz_CtrlState_nextrndKey_428);
    _zz_CtrlState_nextrndKey_429[0] = ((_zz_CtrlState_nextrndKey_425[1] && _zz_CtrlState_nextrndKey_424[1]) ^ _zz_CtrlState_nextrndKey_428);
  end

  assign _zz_CtrlState_nextrndKey_430 = (_zz_CtrlState_nextrndKey_427 ^ _zz_CtrlState_nextrndKey_429);
  always @(*) begin
    _zz_CtrlState_nextrndKey_432[1] = _zz_CtrlState_nextrndKey_430[0];
    _zz_CtrlState_nextrndKey_432[0] = _zz_CtrlState_nextrndKey_430[1];
  end

  assign _zz_CtrlState_nextrndKey_431 = _zz_CtrlState_nextrndKey_432;
  assign _zz_CtrlState_nextrndKey_433 = ((_zz_CtrlState_nextrndKey_431[0] && _zz_CtrlState_nextrndKey_424[1]) ^ (_zz_CtrlState_nextrndKey_424[0] && _zz_CtrlState_nextrndKey_431[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_434[1] = ((_zz_CtrlState_nextrndKey_431[0] && _zz_CtrlState_nextrndKey_424[0]) ^ _zz_CtrlState_nextrndKey_433);
    _zz_CtrlState_nextrndKey_434[0] = ((_zz_CtrlState_nextrndKey_431[1] && _zz_CtrlState_nextrndKey_424[1]) ^ _zz_CtrlState_nextrndKey_433);
  end

  assign _zz_CtrlState_nextrndKey_435 = ((_zz_CtrlState_nextrndKey_431[0] && _zz_CtrlState_nextrndKey_425[1]) ^ (_zz_CtrlState_nextrndKey_425[0] && _zz_CtrlState_nextrndKey_431[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_436[1] = ((_zz_CtrlState_nextrndKey_431[0] && _zz_CtrlState_nextrndKey_425[0]) ^ _zz_CtrlState_nextrndKey_435);
    _zz_CtrlState_nextrndKey_436[0] = ((_zz_CtrlState_nextrndKey_431[1] && _zz_CtrlState_nextrndKey_425[1]) ^ _zz_CtrlState_nextrndKey_435);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_423[3 : 2] = _zz_CtrlState_nextrndKey_436;
    _zz_CtrlState_nextrndKey_423[1 : 0] = _zz_CtrlState_nextrndKey_434;
  end

  assign _zz_CtrlState_nextrndKey_422 = _zz_CtrlState_nextrndKey_423;
  assign _zz_CtrlState_nextrndKey_438 = _zz_CtrlState_nextrndKey_401[3 : 2];
  assign _zz_CtrlState_nextrndKey_439 = _zz_CtrlState_nextrndKey_401[1 : 0];
  assign _zz_CtrlState_nextrndKey_440 = _zz_CtrlState_nextrndKey_422[3 : 2];
  assign _zz_CtrlState_nextrndKey_441 = _zz_CtrlState_nextrndKey_422[1 : 0];
  assign _zz_CtrlState_nextrndKey_442 = (_zz_CtrlState_nextrndKey_438 ^ _zz_CtrlState_nextrndKey_439);
  assign _zz_CtrlState_nextrndKey_443 = (_zz_CtrlState_nextrndKey_440 ^ _zz_CtrlState_nextrndKey_441);
  assign _zz_CtrlState_nextrndKey_445 = ((_zz_CtrlState_nextrndKey_443[0] && _zz_CtrlState_nextrndKey_442[1]) ^ (_zz_CtrlState_nextrndKey_442[0] && _zz_CtrlState_nextrndKey_443[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_446[1] = ((_zz_CtrlState_nextrndKey_443[0] && _zz_CtrlState_nextrndKey_442[0]) ^ _zz_CtrlState_nextrndKey_445);
    _zz_CtrlState_nextrndKey_446[0] = ((_zz_CtrlState_nextrndKey_443[1] && _zz_CtrlState_nextrndKey_442[1]) ^ _zz_CtrlState_nextrndKey_445);
  end

  assign _zz_CtrlState_nextrndKey_444 = _zz_CtrlState_nextrndKey_446;
  always @(*) begin
    _zz_CtrlState_nextrndKey_448[1] = _zz_CtrlState_nextrndKey_444[0];
    _zz_CtrlState_nextrndKey_448[0] = (_zz_CtrlState_nextrndKey_444[0] ^ _zz_CtrlState_nextrndKey_444[1]);
  end

  assign _zz_CtrlState_nextrndKey_447 = _zz_CtrlState_nextrndKey_448;
  assign _zz_CtrlState_nextrndKey_449 = ((_zz_CtrlState_nextrndKey_440[0] && _zz_CtrlState_nextrndKey_438[1]) ^ (_zz_CtrlState_nextrndKey_438[0] && _zz_CtrlState_nextrndKey_440[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_450[1] = ((_zz_CtrlState_nextrndKey_440[0] && _zz_CtrlState_nextrndKey_438[0]) ^ _zz_CtrlState_nextrndKey_449);
    _zz_CtrlState_nextrndKey_450[0] = ((_zz_CtrlState_nextrndKey_440[1] && _zz_CtrlState_nextrndKey_438[1]) ^ _zz_CtrlState_nextrndKey_449);
  end

  assign _zz_CtrlState_nextrndKey_451 = ((_zz_CtrlState_nextrndKey_441[0] && _zz_CtrlState_nextrndKey_439[1]) ^ (_zz_CtrlState_nextrndKey_439[0] && _zz_CtrlState_nextrndKey_441[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_452[1] = ((_zz_CtrlState_nextrndKey_441[0] && _zz_CtrlState_nextrndKey_439[0]) ^ _zz_CtrlState_nextrndKey_451);
    _zz_CtrlState_nextrndKey_452[0] = ((_zz_CtrlState_nextrndKey_441[1] && _zz_CtrlState_nextrndKey_439[1]) ^ _zz_CtrlState_nextrndKey_451);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_437[3 : 2] = (_zz_CtrlState_nextrndKey_450 ^ _zz_CtrlState_nextrndKey_447);
    _zz_CtrlState_nextrndKey_437[1 : 0] = (_zz_CtrlState_nextrndKey_452 ^ _zz_CtrlState_nextrndKey_447);
  end

  assign _zz_CtrlState_nextrndKey_454 = _zz_CtrlState_nextrndKey_402[3 : 2];
  assign _zz_CtrlState_nextrndKey_455 = _zz_CtrlState_nextrndKey_402[1 : 0];
  assign _zz_CtrlState_nextrndKey_456 = _zz_CtrlState_nextrndKey_422[3 : 2];
  assign _zz_CtrlState_nextrndKey_457 = _zz_CtrlState_nextrndKey_422[1 : 0];
  assign _zz_CtrlState_nextrndKey_458 = (_zz_CtrlState_nextrndKey_454 ^ _zz_CtrlState_nextrndKey_455);
  assign _zz_CtrlState_nextrndKey_459 = (_zz_CtrlState_nextrndKey_456 ^ _zz_CtrlState_nextrndKey_457);
  assign _zz_CtrlState_nextrndKey_461 = ((_zz_CtrlState_nextrndKey_459[0] && _zz_CtrlState_nextrndKey_458[1]) ^ (_zz_CtrlState_nextrndKey_458[0] && _zz_CtrlState_nextrndKey_459[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_462[1] = ((_zz_CtrlState_nextrndKey_459[0] && _zz_CtrlState_nextrndKey_458[0]) ^ _zz_CtrlState_nextrndKey_461);
    _zz_CtrlState_nextrndKey_462[0] = ((_zz_CtrlState_nextrndKey_459[1] && _zz_CtrlState_nextrndKey_458[1]) ^ _zz_CtrlState_nextrndKey_461);
  end

  assign _zz_CtrlState_nextrndKey_460 = _zz_CtrlState_nextrndKey_462;
  always @(*) begin
    _zz_CtrlState_nextrndKey_464[1] = _zz_CtrlState_nextrndKey_460[0];
    _zz_CtrlState_nextrndKey_464[0] = (_zz_CtrlState_nextrndKey_460[0] ^ _zz_CtrlState_nextrndKey_460[1]);
  end

  assign _zz_CtrlState_nextrndKey_463 = _zz_CtrlState_nextrndKey_464;
  assign _zz_CtrlState_nextrndKey_465 = ((_zz_CtrlState_nextrndKey_456[0] && _zz_CtrlState_nextrndKey_454[1]) ^ (_zz_CtrlState_nextrndKey_454[0] && _zz_CtrlState_nextrndKey_456[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_466[1] = ((_zz_CtrlState_nextrndKey_456[0] && _zz_CtrlState_nextrndKey_454[0]) ^ _zz_CtrlState_nextrndKey_465);
    _zz_CtrlState_nextrndKey_466[0] = ((_zz_CtrlState_nextrndKey_456[1] && _zz_CtrlState_nextrndKey_454[1]) ^ _zz_CtrlState_nextrndKey_465);
  end

  assign _zz_CtrlState_nextrndKey_467 = ((_zz_CtrlState_nextrndKey_457[0] && _zz_CtrlState_nextrndKey_455[1]) ^ (_zz_CtrlState_nextrndKey_455[0] && _zz_CtrlState_nextrndKey_457[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_468[1] = ((_zz_CtrlState_nextrndKey_457[0] && _zz_CtrlState_nextrndKey_455[0]) ^ _zz_CtrlState_nextrndKey_467);
    _zz_CtrlState_nextrndKey_468[0] = ((_zz_CtrlState_nextrndKey_457[1] && _zz_CtrlState_nextrndKey_455[1]) ^ _zz_CtrlState_nextrndKey_467);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_453[3 : 2] = (_zz_CtrlState_nextrndKey_466 ^ _zz_CtrlState_nextrndKey_463);
    _zz_CtrlState_nextrndKey_453[1 : 0] = (_zz_CtrlState_nextrndKey_468 ^ _zz_CtrlState_nextrndKey_463);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_400[7 : 4] = _zz_CtrlState_nextrndKey_453;
    _zz_CtrlState_nextrndKey_400[3 : 0] = _zz_CtrlState_nextrndKey_437;
  end

  assign _zz_CtrlState_nextrndKey_399 = _zz_CtrlState_nextrndKey_400;
  always @(*) begin
    _zz_CtrlState_nextrndKey_470[7] = (_zz_CtrlState_nextrndKey_399[5] ^ _zz_CtrlState_nextrndKey_399[3]);
    _zz_CtrlState_nextrndKey_470[6] = (_zz_CtrlState_nextrndKey_399[7] ^ _zz_CtrlState_nextrndKey_399[3]);
    _zz_CtrlState_nextrndKey_470[5] = (_zz_CtrlState_nextrndKey_399[6] ^ _zz_CtrlState_nextrndKey_399[0]);
    _zz_CtrlState_nextrndKey_470[4] = ((_zz_CtrlState_nextrndKey_399[7] ^ _zz_CtrlState_nextrndKey_399[5]) ^ _zz_CtrlState_nextrndKey_399[3]);
    _zz_CtrlState_nextrndKey_470[3] = ((((_zz_CtrlState_nextrndKey_399[7] ^ _zz_CtrlState_nextrndKey_399[6]) ^ _zz_CtrlState_nextrndKey_399[5]) ^ _zz_CtrlState_nextrndKey_399[4]) ^ _zz_CtrlState_nextrndKey_399[3]);
    _zz_CtrlState_nextrndKey_470[2] = ((((_zz_CtrlState_nextrndKey_399[6] ^ _zz_CtrlState_nextrndKey_399[5]) ^ _zz_CtrlState_nextrndKey_399[3]) ^ _zz_CtrlState_nextrndKey_399[2]) ^ _zz_CtrlState_nextrndKey_399[0]);
    _zz_CtrlState_nextrndKey_470[1] = ((_zz_CtrlState_nextrndKey_399[5] ^ _zz_CtrlState_nextrndKey_399[4]) ^ _zz_CtrlState_nextrndKey_399[1]);
    _zz_CtrlState_nextrndKey_470[0] = ((_zz_CtrlState_nextrndKey_399[6] ^ _zz_CtrlState_nextrndKey_399[4]) ^ _zz_CtrlState_nextrndKey_399[1]);
  end

  assign _zz_CtrlState_nextrndKey_469 = _zz_CtrlState_nextrndKey_470;
  always @(*) begin
    _zz_CtrlState_nextrndKey_396[7] = _zz_CtrlState_nextrndKey_469[7];
    _zz_CtrlState_nextrndKey_396[6] = (! _zz_CtrlState_nextrndKey_469[6]);
    _zz_CtrlState_nextrndKey_396[5] = (! _zz_CtrlState_nextrndKey_469[5]);
    _zz_CtrlState_nextrndKey_396[4] = _zz_CtrlState_nextrndKey_469[4];
    _zz_CtrlState_nextrndKey_396[3] = _zz_CtrlState_nextrndKey_469[3];
    _zz_CtrlState_nextrndKey_396[2] = _zz_CtrlState_nextrndKey_469[2];
    _zz_CtrlState_nextrndKey_396[1] = (! _zz_CtrlState_nextrndKey_469[1]);
    _zz_CtrlState_nextrndKey_396[0] = (! _zz_CtrlState_nextrndKey_469[0]);
  end

  assign _zz_CtrlState_nextrndKey_471 = _zz_CtrlState_nextrndKey_317[23 : 16];
  always @(*) begin
    _zz_CtrlState_nextrndKey_474[7] = (((((_zz_CtrlState_nextrndKey_471[7] ^ _zz_CtrlState_nextrndKey_471[6]) ^ _zz_CtrlState_nextrndKey_471[5]) ^ _zz_CtrlState_nextrndKey_471[2]) ^ _zz_CtrlState_nextrndKey_471[1]) ^ _zz_CtrlState_nextrndKey_471[0]);
    _zz_CtrlState_nextrndKey_474[6] = (((_zz_CtrlState_nextrndKey_471[6] ^ _zz_CtrlState_nextrndKey_471[5]) ^ _zz_CtrlState_nextrndKey_471[4]) ^ _zz_CtrlState_nextrndKey_471[0]);
    _zz_CtrlState_nextrndKey_474[5] = (((_zz_CtrlState_nextrndKey_471[6] ^ _zz_CtrlState_nextrndKey_471[5]) ^ _zz_CtrlState_nextrndKey_471[1]) ^ _zz_CtrlState_nextrndKey_471[0]);
    _zz_CtrlState_nextrndKey_474[4] = (((_zz_CtrlState_nextrndKey_471[7] ^ _zz_CtrlState_nextrndKey_471[6]) ^ _zz_CtrlState_nextrndKey_471[5]) ^ _zz_CtrlState_nextrndKey_471[0]);
    _zz_CtrlState_nextrndKey_474[3] = ((((_zz_CtrlState_nextrndKey_471[7] ^ _zz_CtrlState_nextrndKey_471[4]) ^ _zz_CtrlState_nextrndKey_471[3]) ^ _zz_CtrlState_nextrndKey_471[1]) ^ _zz_CtrlState_nextrndKey_471[0]);
    _zz_CtrlState_nextrndKey_474[2] = _zz_CtrlState_nextrndKey_471[0];
    _zz_CtrlState_nextrndKey_474[1] = ((_zz_CtrlState_nextrndKey_471[6] ^ _zz_CtrlState_nextrndKey_471[5]) ^ _zz_CtrlState_nextrndKey_471[0]);
    _zz_CtrlState_nextrndKey_474[0] = ((((_zz_CtrlState_nextrndKey_471[6] ^ _zz_CtrlState_nextrndKey_471[3]) ^ _zz_CtrlState_nextrndKey_471[2]) ^ _zz_CtrlState_nextrndKey_471[1]) ^ _zz_CtrlState_nextrndKey_471[0]);
  end

  assign _zz_CtrlState_nextrndKey_473 = _zz_CtrlState_nextrndKey_474;
  assign _zz_CtrlState_nextrndKey_477 = _zz_CtrlState_nextrndKey_473[7 : 4];
  assign _zz_CtrlState_nextrndKey_478 = _zz_CtrlState_nextrndKey_473[3 : 0];
  assign _zz_CtrlState_nextrndKey_479 = (_zz_CtrlState_nextrndKey_477 ^ _zz_CtrlState_nextrndKey_478);
  always @(*) begin
    _zz_CtrlState_nextrndKey_480[3] = (_zz_CtrlState_nextrndKey_479[2] ^ _zz_CtrlState_nextrndKey_479[0]);
    _zz_CtrlState_nextrndKey_480[2] = (_zz_CtrlState_nextrndKey_479[3] ^ _zz_CtrlState_nextrndKey_479[1]);
    _zz_CtrlState_nextrndKey_480[1] = (_zz_CtrlState_nextrndKey_479[1] ^ _zz_CtrlState_nextrndKey_479[0]);
    _zz_CtrlState_nextrndKey_480[0] = _zz_CtrlState_nextrndKey_479[0];
  end

  assign _zz_CtrlState_nextrndKey_482 = _zz_CtrlState_nextrndKey_477[3 : 2];
  assign _zz_CtrlState_nextrndKey_483 = _zz_CtrlState_nextrndKey_477[1 : 0];
  assign _zz_CtrlState_nextrndKey_484 = _zz_CtrlState_nextrndKey_478[3 : 2];
  assign _zz_CtrlState_nextrndKey_485 = _zz_CtrlState_nextrndKey_478[1 : 0];
  assign _zz_CtrlState_nextrndKey_486 = (_zz_CtrlState_nextrndKey_482 ^ _zz_CtrlState_nextrndKey_483);
  assign _zz_CtrlState_nextrndKey_487 = (_zz_CtrlState_nextrndKey_484 ^ _zz_CtrlState_nextrndKey_485);
  assign _zz_CtrlState_nextrndKey_489 = ((_zz_CtrlState_nextrndKey_487[0] && _zz_CtrlState_nextrndKey_486[1]) ^ (_zz_CtrlState_nextrndKey_486[0] && _zz_CtrlState_nextrndKey_487[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_490[1] = ((_zz_CtrlState_nextrndKey_487[0] && _zz_CtrlState_nextrndKey_486[0]) ^ _zz_CtrlState_nextrndKey_489);
    _zz_CtrlState_nextrndKey_490[0] = ((_zz_CtrlState_nextrndKey_487[1] && _zz_CtrlState_nextrndKey_486[1]) ^ _zz_CtrlState_nextrndKey_489);
  end

  assign _zz_CtrlState_nextrndKey_488 = _zz_CtrlState_nextrndKey_490;
  always @(*) begin
    _zz_CtrlState_nextrndKey_492[1] = _zz_CtrlState_nextrndKey_488[0];
    _zz_CtrlState_nextrndKey_492[0] = (_zz_CtrlState_nextrndKey_488[0] ^ _zz_CtrlState_nextrndKey_488[1]);
  end

  assign _zz_CtrlState_nextrndKey_491 = _zz_CtrlState_nextrndKey_492;
  assign _zz_CtrlState_nextrndKey_493 = ((_zz_CtrlState_nextrndKey_484[0] && _zz_CtrlState_nextrndKey_482[1]) ^ (_zz_CtrlState_nextrndKey_482[0] && _zz_CtrlState_nextrndKey_484[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_494[1] = ((_zz_CtrlState_nextrndKey_484[0] && _zz_CtrlState_nextrndKey_482[0]) ^ _zz_CtrlState_nextrndKey_493);
    _zz_CtrlState_nextrndKey_494[0] = ((_zz_CtrlState_nextrndKey_484[1] && _zz_CtrlState_nextrndKey_482[1]) ^ _zz_CtrlState_nextrndKey_493);
  end

  assign _zz_CtrlState_nextrndKey_495 = ((_zz_CtrlState_nextrndKey_485[0] && _zz_CtrlState_nextrndKey_483[1]) ^ (_zz_CtrlState_nextrndKey_483[0] && _zz_CtrlState_nextrndKey_485[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_496[1] = ((_zz_CtrlState_nextrndKey_485[0] && _zz_CtrlState_nextrndKey_483[0]) ^ _zz_CtrlState_nextrndKey_495);
    _zz_CtrlState_nextrndKey_496[0] = ((_zz_CtrlState_nextrndKey_485[1] && _zz_CtrlState_nextrndKey_483[1]) ^ _zz_CtrlState_nextrndKey_495);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_481[3 : 2] = (_zz_CtrlState_nextrndKey_494 ^ _zz_CtrlState_nextrndKey_491);
    _zz_CtrlState_nextrndKey_481[1 : 0] = (_zz_CtrlState_nextrndKey_496 ^ _zz_CtrlState_nextrndKey_491);
  end

  assign _zz_CtrlState_nextrndKey_497 = (_zz_CtrlState_nextrndKey_480 ^ _zz_CtrlState_nextrndKey_481);
  assign _zz_CtrlState_nextrndKey_500 = _zz_CtrlState_nextrndKey_497[3 : 2];
  assign _zz_CtrlState_nextrndKey_501 = _zz_CtrlState_nextrndKey_497[1 : 0];
  assign _zz_CtrlState_nextrndKey_502 = (_zz_CtrlState_nextrndKey_500 ^ _zz_CtrlState_nextrndKey_501);
  always @(*) begin
    _zz_CtrlState_nextrndKey_503[1] = _zz_CtrlState_nextrndKey_502[1];
    _zz_CtrlState_nextrndKey_503[0] = (_zz_CtrlState_nextrndKey_502[0] ^ _zz_CtrlState_nextrndKey_502[1]);
  end

  assign _zz_CtrlState_nextrndKey_504 = ((_zz_CtrlState_nextrndKey_501[0] && _zz_CtrlState_nextrndKey_500[1]) ^ (_zz_CtrlState_nextrndKey_500[0] && _zz_CtrlState_nextrndKey_501[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_505[1] = ((_zz_CtrlState_nextrndKey_501[0] && _zz_CtrlState_nextrndKey_500[0]) ^ _zz_CtrlState_nextrndKey_504);
    _zz_CtrlState_nextrndKey_505[0] = ((_zz_CtrlState_nextrndKey_501[1] && _zz_CtrlState_nextrndKey_500[1]) ^ _zz_CtrlState_nextrndKey_504);
  end

  assign _zz_CtrlState_nextrndKey_506 = (_zz_CtrlState_nextrndKey_503 ^ _zz_CtrlState_nextrndKey_505);
  always @(*) begin
    _zz_CtrlState_nextrndKey_508[1] = _zz_CtrlState_nextrndKey_506[0];
    _zz_CtrlState_nextrndKey_508[0] = _zz_CtrlState_nextrndKey_506[1];
  end

  assign _zz_CtrlState_nextrndKey_507 = _zz_CtrlState_nextrndKey_508;
  assign _zz_CtrlState_nextrndKey_509 = ((_zz_CtrlState_nextrndKey_507[0] && _zz_CtrlState_nextrndKey_500[1]) ^ (_zz_CtrlState_nextrndKey_500[0] && _zz_CtrlState_nextrndKey_507[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_510[1] = ((_zz_CtrlState_nextrndKey_507[0] && _zz_CtrlState_nextrndKey_500[0]) ^ _zz_CtrlState_nextrndKey_509);
    _zz_CtrlState_nextrndKey_510[0] = ((_zz_CtrlState_nextrndKey_507[1] && _zz_CtrlState_nextrndKey_500[1]) ^ _zz_CtrlState_nextrndKey_509);
  end

  assign _zz_CtrlState_nextrndKey_511 = ((_zz_CtrlState_nextrndKey_507[0] && _zz_CtrlState_nextrndKey_501[1]) ^ (_zz_CtrlState_nextrndKey_501[0] && _zz_CtrlState_nextrndKey_507[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_512[1] = ((_zz_CtrlState_nextrndKey_507[0] && _zz_CtrlState_nextrndKey_501[0]) ^ _zz_CtrlState_nextrndKey_511);
    _zz_CtrlState_nextrndKey_512[0] = ((_zz_CtrlState_nextrndKey_507[1] && _zz_CtrlState_nextrndKey_501[1]) ^ _zz_CtrlState_nextrndKey_511);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_499[3 : 2] = _zz_CtrlState_nextrndKey_512;
    _zz_CtrlState_nextrndKey_499[1 : 0] = _zz_CtrlState_nextrndKey_510;
  end

  assign _zz_CtrlState_nextrndKey_498 = _zz_CtrlState_nextrndKey_499;
  assign _zz_CtrlState_nextrndKey_514 = _zz_CtrlState_nextrndKey_477[3 : 2];
  assign _zz_CtrlState_nextrndKey_515 = _zz_CtrlState_nextrndKey_477[1 : 0];
  assign _zz_CtrlState_nextrndKey_516 = _zz_CtrlState_nextrndKey_498[3 : 2];
  assign _zz_CtrlState_nextrndKey_517 = _zz_CtrlState_nextrndKey_498[1 : 0];
  assign _zz_CtrlState_nextrndKey_518 = (_zz_CtrlState_nextrndKey_514 ^ _zz_CtrlState_nextrndKey_515);
  assign _zz_CtrlState_nextrndKey_519 = (_zz_CtrlState_nextrndKey_516 ^ _zz_CtrlState_nextrndKey_517);
  assign _zz_CtrlState_nextrndKey_521 = ((_zz_CtrlState_nextrndKey_519[0] && _zz_CtrlState_nextrndKey_518[1]) ^ (_zz_CtrlState_nextrndKey_518[0] && _zz_CtrlState_nextrndKey_519[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_522[1] = ((_zz_CtrlState_nextrndKey_519[0] && _zz_CtrlState_nextrndKey_518[0]) ^ _zz_CtrlState_nextrndKey_521);
    _zz_CtrlState_nextrndKey_522[0] = ((_zz_CtrlState_nextrndKey_519[1] && _zz_CtrlState_nextrndKey_518[1]) ^ _zz_CtrlState_nextrndKey_521);
  end

  assign _zz_CtrlState_nextrndKey_520 = _zz_CtrlState_nextrndKey_522;
  always @(*) begin
    _zz_CtrlState_nextrndKey_524[1] = _zz_CtrlState_nextrndKey_520[0];
    _zz_CtrlState_nextrndKey_524[0] = (_zz_CtrlState_nextrndKey_520[0] ^ _zz_CtrlState_nextrndKey_520[1]);
  end

  assign _zz_CtrlState_nextrndKey_523 = _zz_CtrlState_nextrndKey_524;
  assign _zz_CtrlState_nextrndKey_525 = ((_zz_CtrlState_nextrndKey_516[0] && _zz_CtrlState_nextrndKey_514[1]) ^ (_zz_CtrlState_nextrndKey_514[0] && _zz_CtrlState_nextrndKey_516[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_526[1] = ((_zz_CtrlState_nextrndKey_516[0] && _zz_CtrlState_nextrndKey_514[0]) ^ _zz_CtrlState_nextrndKey_525);
    _zz_CtrlState_nextrndKey_526[0] = ((_zz_CtrlState_nextrndKey_516[1] && _zz_CtrlState_nextrndKey_514[1]) ^ _zz_CtrlState_nextrndKey_525);
  end

  assign _zz_CtrlState_nextrndKey_527 = ((_zz_CtrlState_nextrndKey_517[0] && _zz_CtrlState_nextrndKey_515[1]) ^ (_zz_CtrlState_nextrndKey_515[0] && _zz_CtrlState_nextrndKey_517[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_528[1] = ((_zz_CtrlState_nextrndKey_517[0] && _zz_CtrlState_nextrndKey_515[0]) ^ _zz_CtrlState_nextrndKey_527);
    _zz_CtrlState_nextrndKey_528[0] = ((_zz_CtrlState_nextrndKey_517[1] && _zz_CtrlState_nextrndKey_515[1]) ^ _zz_CtrlState_nextrndKey_527);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_513[3 : 2] = (_zz_CtrlState_nextrndKey_526 ^ _zz_CtrlState_nextrndKey_523);
    _zz_CtrlState_nextrndKey_513[1 : 0] = (_zz_CtrlState_nextrndKey_528 ^ _zz_CtrlState_nextrndKey_523);
  end

  assign _zz_CtrlState_nextrndKey_530 = _zz_CtrlState_nextrndKey_478[3 : 2];
  assign _zz_CtrlState_nextrndKey_531 = _zz_CtrlState_nextrndKey_478[1 : 0];
  assign _zz_CtrlState_nextrndKey_532 = _zz_CtrlState_nextrndKey_498[3 : 2];
  assign _zz_CtrlState_nextrndKey_533 = _zz_CtrlState_nextrndKey_498[1 : 0];
  assign _zz_CtrlState_nextrndKey_534 = (_zz_CtrlState_nextrndKey_530 ^ _zz_CtrlState_nextrndKey_531);
  assign _zz_CtrlState_nextrndKey_535 = (_zz_CtrlState_nextrndKey_532 ^ _zz_CtrlState_nextrndKey_533);
  assign _zz_CtrlState_nextrndKey_537 = ((_zz_CtrlState_nextrndKey_535[0] && _zz_CtrlState_nextrndKey_534[1]) ^ (_zz_CtrlState_nextrndKey_534[0] && _zz_CtrlState_nextrndKey_535[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_538[1] = ((_zz_CtrlState_nextrndKey_535[0] && _zz_CtrlState_nextrndKey_534[0]) ^ _zz_CtrlState_nextrndKey_537);
    _zz_CtrlState_nextrndKey_538[0] = ((_zz_CtrlState_nextrndKey_535[1] && _zz_CtrlState_nextrndKey_534[1]) ^ _zz_CtrlState_nextrndKey_537);
  end

  assign _zz_CtrlState_nextrndKey_536 = _zz_CtrlState_nextrndKey_538;
  always @(*) begin
    _zz_CtrlState_nextrndKey_540[1] = _zz_CtrlState_nextrndKey_536[0];
    _zz_CtrlState_nextrndKey_540[0] = (_zz_CtrlState_nextrndKey_536[0] ^ _zz_CtrlState_nextrndKey_536[1]);
  end

  assign _zz_CtrlState_nextrndKey_539 = _zz_CtrlState_nextrndKey_540;
  assign _zz_CtrlState_nextrndKey_541 = ((_zz_CtrlState_nextrndKey_532[0] && _zz_CtrlState_nextrndKey_530[1]) ^ (_zz_CtrlState_nextrndKey_530[0] && _zz_CtrlState_nextrndKey_532[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_542[1] = ((_zz_CtrlState_nextrndKey_532[0] && _zz_CtrlState_nextrndKey_530[0]) ^ _zz_CtrlState_nextrndKey_541);
    _zz_CtrlState_nextrndKey_542[0] = ((_zz_CtrlState_nextrndKey_532[1] && _zz_CtrlState_nextrndKey_530[1]) ^ _zz_CtrlState_nextrndKey_541);
  end

  assign _zz_CtrlState_nextrndKey_543 = ((_zz_CtrlState_nextrndKey_533[0] && _zz_CtrlState_nextrndKey_531[1]) ^ (_zz_CtrlState_nextrndKey_531[0] && _zz_CtrlState_nextrndKey_533[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_544[1] = ((_zz_CtrlState_nextrndKey_533[0] && _zz_CtrlState_nextrndKey_531[0]) ^ _zz_CtrlState_nextrndKey_543);
    _zz_CtrlState_nextrndKey_544[0] = ((_zz_CtrlState_nextrndKey_533[1] && _zz_CtrlState_nextrndKey_531[1]) ^ _zz_CtrlState_nextrndKey_543);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_529[3 : 2] = (_zz_CtrlState_nextrndKey_542 ^ _zz_CtrlState_nextrndKey_539);
    _zz_CtrlState_nextrndKey_529[1 : 0] = (_zz_CtrlState_nextrndKey_544 ^ _zz_CtrlState_nextrndKey_539);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_476[7 : 4] = _zz_CtrlState_nextrndKey_529;
    _zz_CtrlState_nextrndKey_476[3 : 0] = _zz_CtrlState_nextrndKey_513;
  end

  assign _zz_CtrlState_nextrndKey_475 = _zz_CtrlState_nextrndKey_476;
  always @(*) begin
    _zz_CtrlState_nextrndKey_546[7] = (_zz_CtrlState_nextrndKey_475[5] ^ _zz_CtrlState_nextrndKey_475[3]);
    _zz_CtrlState_nextrndKey_546[6] = (_zz_CtrlState_nextrndKey_475[7] ^ _zz_CtrlState_nextrndKey_475[3]);
    _zz_CtrlState_nextrndKey_546[5] = (_zz_CtrlState_nextrndKey_475[6] ^ _zz_CtrlState_nextrndKey_475[0]);
    _zz_CtrlState_nextrndKey_546[4] = ((_zz_CtrlState_nextrndKey_475[7] ^ _zz_CtrlState_nextrndKey_475[5]) ^ _zz_CtrlState_nextrndKey_475[3]);
    _zz_CtrlState_nextrndKey_546[3] = ((((_zz_CtrlState_nextrndKey_475[7] ^ _zz_CtrlState_nextrndKey_475[6]) ^ _zz_CtrlState_nextrndKey_475[5]) ^ _zz_CtrlState_nextrndKey_475[4]) ^ _zz_CtrlState_nextrndKey_475[3]);
    _zz_CtrlState_nextrndKey_546[2] = ((((_zz_CtrlState_nextrndKey_475[6] ^ _zz_CtrlState_nextrndKey_475[5]) ^ _zz_CtrlState_nextrndKey_475[3]) ^ _zz_CtrlState_nextrndKey_475[2]) ^ _zz_CtrlState_nextrndKey_475[0]);
    _zz_CtrlState_nextrndKey_546[1] = ((_zz_CtrlState_nextrndKey_475[5] ^ _zz_CtrlState_nextrndKey_475[4]) ^ _zz_CtrlState_nextrndKey_475[1]);
    _zz_CtrlState_nextrndKey_546[0] = ((_zz_CtrlState_nextrndKey_475[6] ^ _zz_CtrlState_nextrndKey_475[4]) ^ _zz_CtrlState_nextrndKey_475[1]);
  end

  assign _zz_CtrlState_nextrndKey_545 = _zz_CtrlState_nextrndKey_546;
  always @(*) begin
    _zz_CtrlState_nextrndKey_472[7] = _zz_CtrlState_nextrndKey_545[7];
    _zz_CtrlState_nextrndKey_472[6] = (! _zz_CtrlState_nextrndKey_545[6]);
    _zz_CtrlState_nextrndKey_472[5] = (! _zz_CtrlState_nextrndKey_545[5]);
    _zz_CtrlState_nextrndKey_472[4] = _zz_CtrlState_nextrndKey_545[4];
    _zz_CtrlState_nextrndKey_472[3] = _zz_CtrlState_nextrndKey_545[3];
    _zz_CtrlState_nextrndKey_472[2] = _zz_CtrlState_nextrndKey_545[2];
    _zz_CtrlState_nextrndKey_472[1] = (! _zz_CtrlState_nextrndKey_545[1]);
    _zz_CtrlState_nextrndKey_472[0] = (! _zz_CtrlState_nextrndKey_545[0]);
  end

  assign _zz_CtrlState_nextrndKey_547 = _zz_CtrlState_nextrndKey_317[31 : 24];
  always @(*) begin
    _zz_CtrlState_nextrndKey_550[7] = (((((_zz_CtrlState_nextrndKey_547[7] ^ _zz_CtrlState_nextrndKey_547[6]) ^ _zz_CtrlState_nextrndKey_547[5]) ^ _zz_CtrlState_nextrndKey_547[2]) ^ _zz_CtrlState_nextrndKey_547[1]) ^ _zz_CtrlState_nextrndKey_547[0]);
    _zz_CtrlState_nextrndKey_550[6] = (((_zz_CtrlState_nextrndKey_547[6] ^ _zz_CtrlState_nextrndKey_547[5]) ^ _zz_CtrlState_nextrndKey_547[4]) ^ _zz_CtrlState_nextrndKey_547[0]);
    _zz_CtrlState_nextrndKey_550[5] = (((_zz_CtrlState_nextrndKey_547[6] ^ _zz_CtrlState_nextrndKey_547[5]) ^ _zz_CtrlState_nextrndKey_547[1]) ^ _zz_CtrlState_nextrndKey_547[0]);
    _zz_CtrlState_nextrndKey_550[4] = (((_zz_CtrlState_nextrndKey_547[7] ^ _zz_CtrlState_nextrndKey_547[6]) ^ _zz_CtrlState_nextrndKey_547[5]) ^ _zz_CtrlState_nextrndKey_547[0]);
    _zz_CtrlState_nextrndKey_550[3] = ((((_zz_CtrlState_nextrndKey_547[7] ^ _zz_CtrlState_nextrndKey_547[4]) ^ _zz_CtrlState_nextrndKey_547[3]) ^ _zz_CtrlState_nextrndKey_547[1]) ^ _zz_CtrlState_nextrndKey_547[0]);
    _zz_CtrlState_nextrndKey_550[2] = _zz_CtrlState_nextrndKey_547[0];
    _zz_CtrlState_nextrndKey_550[1] = ((_zz_CtrlState_nextrndKey_547[6] ^ _zz_CtrlState_nextrndKey_547[5]) ^ _zz_CtrlState_nextrndKey_547[0]);
    _zz_CtrlState_nextrndKey_550[0] = ((((_zz_CtrlState_nextrndKey_547[6] ^ _zz_CtrlState_nextrndKey_547[3]) ^ _zz_CtrlState_nextrndKey_547[2]) ^ _zz_CtrlState_nextrndKey_547[1]) ^ _zz_CtrlState_nextrndKey_547[0]);
  end

  assign _zz_CtrlState_nextrndKey_549 = _zz_CtrlState_nextrndKey_550;
  assign _zz_CtrlState_nextrndKey_553 = _zz_CtrlState_nextrndKey_549[7 : 4];
  assign _zz_CtrlState_nextrndKey_554 = _zz_CtrlState_nextrndKey_549[3 : 0];
  assign _zz_CtrlState_nextrndKey_555 = (_zz_CtrlState_nextrndKey_553 ^ _zz_CtrlState_nextrndKey_554);
  always @(*) begin
    _zz_CtrlState_nextrndKey_556[3] = (_zz_CtrlState_nextrndKey_555[2] ^ _zz_CtrlState_nextrndKey_555[0]);
    _zz_CtrlState_nextrndKey_556[2] = (_zz_CtrlState_nextrndKey_555[3] ^ _zz_CtrlState_nextrndKey_555[1]);
    _zz_CtrlState_nextrndKey_556[1] = (_zz_CtrlState_nextrndKey_555[1] ^ _zz_CtrlState_nextrndKey_555[0]);
    _zz_CtrlState_nextrndKey_556[0] = _zz_CtrlState_nextrndKey_555[0];
  end

  assign _zz_CtrlState_nextrndKey_558 = _zz_CtrlState_nextrndKey_553[3 : 2];
  assign _zz_CtrlState_nextrndKey_559 = _zz_CtrlState_nextrndKey_553[1 : 0];
  assign _zz_CtrlState_nextrndKey_560 = _zz_CtrlState_nextrndKey_554[3 : 2];
  assign _zz_CtrlState_nextrndKey_561 = _zz_CtrlState_nextrndKey_554[1 : 0];
  assign _zz_CtrlState_nextrndKey_562 = (_zz_CtrlState_nextrndKey_558 ^ _zz_CtrlState_nextrndKey_559);
  assign _zz_CtrlState_nextrndKey_563 = (_zz_CtrlState_nextrndKey_560 ^ _zz_CtrlState_nextrndKey_561);
  assign _zz_CtrlState_nextrndKey_565 = ((_zz_CtrlState_nextrndKey_563[0] && _zz_CtrlState_nextrndKey_562[1]) ^ (_zz_CtrlState_nextrndKey_562[0] && _zz_CtrlState_nextrndKey_563[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_566[1] = ((_zz_CtrlState_nextrndKey_563[0] && _zz_CtrlState_nextrndKey_562[0]) ^ _zz_CtrlState_nextrndKey_565);
    _zz_CtrlState_nextrndKey_566[0] = ((_zz_CtrlState_nextrndKey_563[1] && _zz_CtrlState_nextrndKey_562[1]) ^ _zz_CtrlState_nextrndKey_565);
  end

  assign _zz_CtrlState_nextrndKey_564 = _zz_CtrlState_nextrndKey_566;
  always @(*) begin
    _zz_CtrlState_nextrndKey_568[1] = _zz_CtrlState_nextrndKey_564[0];
    _zz_CtrlState_nextrndKey_568[0] = (_zz_CtrlState_nextrndKey_564[0] ^ _zz_CtrlState_nextrndKey_564[1]);
  end

  assign _zz_CtrlState_nextrndKey_567 = _zz_CtrlState_nextrndKey_568;
  assign _zz_CtrlState_nextrndKey_569 = ((_zz_CtrlState_nextrndKey_560[0] && _zz_CtrlState_nextrndKey_558[1]) ^ (_zz_CtrlState_nextrndKey_558[0] && _zz_CtrlState_nextrndKey_560[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_570[1] = ((_zz_CtrlState_nextrndKey_560[0] && _zz_CtrlState_nextrndKey_558[0]) ^ _zz_CtrlState_nextrndKey_569);
    _zz_CtrlState_nextrndKey_570[0] = ((_zz_CtrlState_nextrndKey_560[1] && _zz_CtrlState_nextrndKey_558[1]) ^ _zz_CtrlState_nextrndKey_569);
  end

  assign _zz_CtrlState_nextrndKey_571 = ((_zz_CtrlState_nextrndKey_561[0] && _zz_CtrlState_nextrndKey_559[1]) ^ (_zz_CtrlState_nextrndKey_559[0] && _zz_CtrlState_nextrndKey_561[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_572[1] = ((_zz_CtrlState_nextrndKey_561[0] && _zz_CtrlState_nextrndKey_559[0]) ^ _zz_CtrlState_nextrndKey_571);
    _zz_CtrlState_nextrndKey_572[0] = ((_zz_CtrlState_nextrndKey_561[1] && _zz_CtrlState_nextrndKey_559[1]) ^ _zz_CtrlState_nextrndKey_571);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_557[3 : 2] = (_zz_CtrlState_nextrndKey_570 ^ _zz_CtrlState_nextrndKey_567);
    _zz_CtrlState_nextrndKey_557[1 : 0] = (_zz_CtrlState_nextrndKey_572 ^ _zz_CtrlState_nextrndKey_567);
  end

  assign _zz_CtrlState_nextrndKey_573 = (_zz_CtrlState_nextrndKey_556 ^ _zz_CtrlState_nextrndKey_557);
  assign _zz_CtrlState_nextrndKey_576 = _zz_CtrlState_nextrndKey_573[3 : 2];
  assign _zz_CtrlState_nextrndKey_577 = _zz_CtrlState_nextrndKey_573[1 : 0];
  assign _zz_CtrlState_nextrndKey_578 = (_zz_CtrlState_nextrndKey_576 ^ _zz_CtrlState_nextrndKey_577);
  always @(*) begin
    _zz_CtrlState_nextrndKey_579[1] = _zz_CtrlState_nextrndKey_578[1];
    _zz_CtrlState_nextrndKey_579[0] = (_zz_CtrlState_nextrndKey_578[0] ^ _zz_CtrlState_nextrndKey_578[1]);
  end

  assign _zz_CtrlState_nextrndKey_580 = ((_zz_CtrlState_nextrndKey_577[0] && _zz_CtrlState_nextrndKey_576[1]) ^ (_zz_CtrlState_nextrndKey_576[0] && _zz_CtrlState_nextrndKey_577[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_581[1] = ((_zz_CtrlState_nextrndKey_577[0] && _zz_CtrlState_nextrndKey_576[0]) ^ _zz_CtrlState_nextrndKey_580);
    _zz_CtrlState_nextrndKey_581[0] = ((_zz_CtrlState_nextrndKey_577[1] && _zz_CtrlState_nextrndKey_576[1]) ^ _zz_CtrlState_nextrndKey_580);
  end

  assign _zz_CtrlState_nextrndKey_582 = (_zz_CtrlState_nextrndKey_579 ^ _zz_CtrlState_nextrndKey_581);
  always @(*) begin
    _zz_CtrlState_nextrndKey_584[1] = _zz_CtrlState_nextrndKey_582[0];
    _zz_CtrlState_nextrndKey_584[0] = _zz_CtrlState_nextrndKey_582[1];
  end

  assign _zz_CtrlState_nextrndKey_583 = _zz_CtrlState_nextrndKey_584;
  assign _zz_CtrlState_nextrndKey_585 = ((_zz_CtrlState_nextrndKey_583[0] && _zz_CtrlState_nextrndKey_576[1]) ^ (_zz_CtrlState_nextrndKey_576[0] && _zz_CtrlState_nextrndKey_583[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_586[1] = ((_zz_CtrlState_nextrndKey_583[0] && _zz_CtrlState_nextrndKey_576[0]) ^ _zz_CtrlState_nextrndKey_585);
    _zz_CtrlState_nextrndKey_586[0] = ((_zz_CtrlState_nextrndKey_583[1] && _zz_CtrlState_nextrndKey_576[1]) ^ _zz_CtrlState_nextrndKey_585);
  end

  assign _zz_CtrlState_nextrndKey_587 = ((_zz_CtrlState_nextrndKey_583[0] && _zz_CtrlState_nextrndKey_577[1]) ^ (_zz_CtrlState_nextrndKey_577[0] && _zz_CtrlState_nextrndKey_583[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_588[1] = ((_zz_CtrlState_nextrndKey_583[0] && _zz_CtrlState_nextrndKey_577[0]) ^ _zz_CtrlState_nextrndKey_587);
    _zz_CtrlState_nextrndKey_588[0] = ((_zz_CtrlState_nextrndKey_583[1] && _zz_CtrlState_nextrndKey_577[1]) ^ _zz_CtrlState_nextrndKey_587);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_575[3 : 2] = _zz_CtrlState_nextrndKey_588;
    _zz_CtrlState_nextrndKey_575[1 : 0] = _zz_CtrlState_nextrndKey_586;
  end

  assign _zz_CtrlState_nextrndKey_574 = _zz_CtrlState_nextrndKey_575;
  assign _zz_CtrlState_nextrndKey_590 = _zz_CtrlState_nextrndKey_553[3 : 2];
  assign _zz_CtrlState_nextrndKey_591 = _zz_CtrlState_nextrndKey_553[1 : 0];
  assign _zz_CtrlState_nextrndKey_592 = _zz_CtrlState_nextrndKey_574[3 : 2];
  assign _zz_CtrlState_nextrndKey_593 = _zz_CtrlState_nextrndKey_574[1 : 0];
  assign _zz_CtrlState_nextrndKey_594 = (_zz_CtrlState_nextrndKey_590 ^ _zz_CtrlState_nextrndKey_591);
  assign _zz_CtrlState_nextrndKey_595 = (_zz_CtrlState_nextrndKey_592 ^ _zz_CtrlState_nextrndKey_593);
  assign _zz_CtrlState_nextrndKey_597 = ((_zz_CtrlState_nextrndKey_595[0] && _zz_CtrlState_nextrndKey_594[1]) ^ (_zz_CtrlState_nextrndKey_594[0] && _zz_CtrlState_nextrndKey_595[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_598[1] = ((_zz_CtrlState_nextrndKey_595[0] && _zz_CtrlState_nextrndKey_594[0]) ^ _zz_CtrlState_nextrndKey_597);
    _zz_CtrlState_nextrndKey_598[0] = ((_zz_CtrlState_nextrndKey_595[1] && _zz_CtrlState_nextrndKey_594[1]) ^ _zz_CtrlState_nextrndKey_597);
  end

  assign _zz_CtrlState_nextrndKey_596 = _zz_CtrlState_nextrndKey_598;
  always @(*) begin
    _zz_CtrlState_nextrndKey_600[1] = _zz_CtrlState_nextrndKey_596[0];
    _zz_CtrlState_nextrndKey_600[0] = (_zz_CtrlState_nextrndKey_596[0] ^ _zz_CtrlState_nextrndKey_596[1]);
  end

  assign _zz_CtrlState_nextrndKey_599 = _zz_CtrlState_nextrndKey_600;
  assign _zz_CtrlState_nextrndKey_601 = ((_zz_CtrlState_nextrndKey_592[0] && _zz_CtrlState_nextrndKey_590[1]) ^ (_zz_CtrlState_nextrndKey_590[0] && _zz_CtrlState_nextrndKey_592[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_602[1] = ((_zz_CtrlState_nextrndKey_592[0] && _zz_CtrlState_nextrndKey_590[0]) ^ _zz_CtrlState_nextrndKey_601);
    _zz_CtrlState_nextrndKey_602[0] = ((_zz_CtrlState_nextrndKey_592[1] && _zz_CtrlState_nextrndKey_590[1]) ^ _zz_CtrlState_nextrndKey_601);
  end

  assign _zz_CtrlState_nextrndKey_603 = ((_zz_CtrlState_nextrndKey_593[0] && _zz_CtrlState_nextrndKey_591[1]) ^ (_zz_CtrlState_nextrndKey_591[0] && _zz_CtrlState_nextrndKey_593[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_604[1] = ((_zz_CtrlState_nextrndKey_593[0] && _zz_CtrlState_nextrndKey_591[0]) ^ _zz_CtrlState_nextrndKey_603);
    _zz_CtrlState_nextrndKey_604[0] = ((_zz_CtrlState_nextrndKey_593[1] && _zz_CtrlState_nextrndKey_591[1]) ^ _zz_CtrlState_nextrndKey_603);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_589[3 : 2] = (_zz_CtrlState_nextrndKey_602 ^ _zz_CtrlState_nextrndKey_599);
    _zz_CtrlState_nextrndKey_589[1 : 0] = (_zz_CtrlState_nextrndKey_604 ^ _zz_CtrlState_nextrndKey_599);
  end

  assign _zz_CtrlState_nextrndKey_606 = _zz_CtrlState_nextrndKey_554[3 : 2];
  assign _zz_CtrlState_nextrndKey_607 = _zz_CtrlState_nextrndKey_554[1 : 0];
  assign _zz_CtrlState_nextrndKey_608 = _zz_CtrlState_nextrndKey_574[3 : 2];
  assign _zz_CtrlState_nextrndKey_609 = _zz_CtrlState_nextrndKey_574[1 : 0];
  assign _zz_CtrlState_nextrndKey_610 = (_zz_CtrlState_nextrndKey_606 ^ _zz_CtrlState_nextrndKey_607);
  assign _zz_CtrlState_nextrndKey_611 = (_zz_CtrlState_nextrndKey_608 ^ _zz_CtrlState_nextrndKey_609);
  assign _zz_CtrlState_nextrndKey_613 = ((_zz_CtrlState_nextrndKey_611[0] && _zz_CtrlState_nextrndKey_610[1]) ^ (_zz_CtrlState_nextrndKey_610[0] && _zz_CtrlState_nextrndKey_611[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_614[1] = ((_zz_CtrlState_nextrndKey_611[0] && _zz_CtrlState_nextrndKey_610[0]) ^ _zz_CtrlState_nextrndKey_613);
    _zz_CtrlState_nextrndKey_614[0] = ((_zz_CtrlState_nextrndKey_611[1] && _zz_CtrlState_nextrndKey_610[1]) ^ _zz_CtrlState_nextrndKey_613);
  end

  assign _zz_CtrlState_nextrndKey_612 = _zz_CtrlState_nextrndKey_614;
  always @(*) begin
    _zz_CtrlState_nextrndKey_616[1] = _zz_CtrlState_nextrndKey_612[0];
    _zz_CtrlState_nextrndKey_616[0] = (_zz_CtrlState_nextrndKey_612[0] ^ _zz_CtrlState_nextrndKey_612[1]);
  end

  assign _zz_CtrlState_nextrndKey_615 = _zz_CtrlState_nextrndKey_616;
  assign _zz_CtrlState_nextrndKey_617 = ((_zz_CtrlState_nextrndKey_608[0] && _zz_CtrlState_nextrndKey_606[1]) ^ (_zz_CtrlState_nextrndKey_606[0] && _zz_CtrlState_nextrndKey_608[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_618[1] = ((_zz_CtrlState_nextrndKey_608[0] && _zz_CtrlState_nextrndKey_606[0]) ^ _zz_CtrlState_nextrndKey_617);
    _zz_CtrlState_nextrndKey_618[0] = ((_zz_CtrlState_nextrndKey_608[1] && _zz_CtrlState_nextrndKey_606[1]) ^ _zz_CtrlState_nextrndKey_617);
  end

  assign _zz_CtrlState_nextrndKey_619 = ((_zz_CtrlState_nextrndKey_609[0] && _zz_CtrlState_nextrndKey_607[1]) ^ (_zz_CtrlState_nextrndKey_607[0] && _zz_CtrlState_nextrndKey_609[1]));
  always @(*) begin
    _zz_CtrlState_nextrndKey_620[1] = ((_zz_CtrlState_nextrndKey_609[0] && _zz_CtrlState_nextrndKey_607[0]) ^ _zz_CtrlState_nextrndKey_619);
    _zz_CtrlState_nextrndKey_620[0] = ((_zz_CtrlState_nextrndKey_609[1] && _zz_CtrlState_nextrndKey_607[1]) ^ _zz_CtrlState_nextrndKey_619);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_605[3 : 2] = (_zz_CtrlState_nextrndKey_618 ^ _zz_CtrlState_nextrndKey_615);
    _zz_CtrlState_nextrndKey_605[1 : 0] = (_zz_CtrlState_nextrndKey_620 ^ _zz_CtrlState_nextrndKey_615);
  end

  always @(*) begin
    _zz_CtrlState_nextrndKey_552[7 : 4] = _zz_CtrlState_nextrndKey_605;
    _zz_CtrlState_nextrndKey_552[3 : 0] = _zz_CtrlState_nextrndKey_589;
  end

  assign _zz_CtrlState_nextrndKey_551 = _zz_CtrlState_nextrndKey_552;
  always @(*) begin
    _zz_CtrlState_nextrndKey_622[7] = (_zz_CtrlState_nextrndKey_551[5] ^ _zz_CtrlState_nextrndKey_551[3]);
    _zz_CtrlState_nextrndKey_622[6] = (_zz_CtrlState_nextrndKey_551[7] ^ _zz_CtrlState_nextrndKey_551[3]);
    _zz_CtrlState_nextrndKey_622[5] = (_zz_CtrlState_nextrndKey_551[6] ^ _zz_CtrlState_nextrndKey_551[0]);
    _zz_CtrlState_nextrndKey_622[4] = ((_zz_CtrlState_nextrndKey_551[7] ^ _zz_CtrlState_nextrndKey_551[5]) ^ _zz_CtrlState_nextrndKey_551[3]);
    _zz_CtrlState_nextrndKey_622[3] = ((((_zz_CtrlState_nextrndKey_551[7] ^ _zz_CtrlState_nextrndKey_551[6]) ^ _zz_CtrlState_nextrndKey_551[5]) ^ _zz_CtrlState_nextrndKey_551[4]) ^ _zz_CtrlState_nextrndKey_551[3]);
    _zz_CtrlState_nextrndKey_622[2] = ((((_zz_CtrlState_nextrndKey_551[6] ^ _zz_CtrlState_nextrndKey_551[5]) ^ _zz_CtrlState_nextrndKey_551[3]) ^ _zz_CtrlState_nextrndKey_551[2]) ^ _zz_CtrlState_nextrndKey_551[0]);
    _zz_CtrlState_nextrndKey_622[1] = ((_zz_CtrlState_nextrndKey_551[5] ^ _zz_CtrlState_nextrndKey_551[4]) ^ _zz_CtrlState_nextrndKey_551[1]);
    _zz_CtrlState_nextrndKey_622[0] = ((_zz_CtrlState_nextrndKey_551[6] ^ _zz_CtrlState_nextrndKey_551[4]) ^ _zz_CtrlState_nextrndKey_551[1]);
  end

  assign _zz_CtrlState_nextrndKey_621 = _zz_CtrlState_nextrndKey_622;
  always @(*) begin
    _zz_CtrlState_nextrndKey_548[7] = _zz_CtrlState_nextrndKey_621[7];
    _zz_CtrlState_nextrndKey_548[6] = (! _zz_CtrlState_nextrndKey_621[6]);
    _zz_CtrlState_nextrndKey_548[5] = (! _zz_CtrlState_nextrndKey_621[5]);
    _zz_CtrlState_nextrndKey_548[4] = _zz_CtrlState_nextrndKey_621[4];
    _zz_CtrlState_nextrndKey_548[3] = _zz_CtrlState_nextrndKey_621[3];
    _zz_CtrlState_nextrndKey_548[2] = _zz_CtrlState_nextrndKey_621[2];
    _zz_CtrlState_nextrndKey_548[1] = (! _zz_CtrlState_nextrndKey_621[1]);
    _zz_CtrlState_nextrndKey_548[0] = (! _zz_CtrlState_nextrndKey_621[0]);
  end

  assign _zz_CtrlState_nextrndKey_313 = (_zz_CtrlState_nextrndKey_311[31 : 0] ^ {(_zz_CtrlState_nextrndKey_318[31 : 24] ^ _zz_CtrlState_keyRcon_port0),{_zz_CtrlState_nextrndKey_318[23 : 16],{_zz_CtrlState_nextrndKey_318[15 : 8],_zz_CtrlState_nextrndKey_318[7 : 0]}}});
  assign _zz_CtrlState_nextrndKey_314 = (_zz_CtrlState_nextrndKey_311[63 : 32] ^ _zz_CtrlState_nextrndKey_313);
  assign _zz_CtrlState_nextrndKey_315 = (_zz_CtrlState_nextrndKey_311[95 : 64] ^ _zz_CtrlState_nextrndKey_314);
  assign when_AES_CORE_l78 = (! CtrlState_lastRound);
  assign io_engine_cmd_ready = CtrlState_enginRdy;
  assign io_engine_rsp_payload_block = (CtrlState_dataBuf ^ CtrlState_nextrndKey);
  assign io_engine_rsp_valid = CtrlState_lastRound_regNext;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      CtrlState_enginRdy <= 1'b1;
      CtrlState_ongoing <= 1'b0;
      CtrlState_nextrndKey <= 128'h0;
      CtrlState_rndCnt <= 4'b0000;
      CtrlState_dataBuf <= 128'h0;
      CtrlState_lastRound_regNext <= 1'b0;
    end else begin
      if(io_engine_cmd_fire_1) begin
        CtrlState_ongoing <= 1'b1;
        CtrlState_enginRdy <= 1'b0;
        CtrlState_rndCnt <= 4'b0001;
        CtrlState_nextrndKey <= {_zz_CtrlState_nextrndKey_1,{_zz_CtrlState_nextrndKey_2,{_zz_CtrlState_nextrndKey_3,(_zz_CtrlState_nextrndKey_4 ^ _zz_CtrlState_nextrndKey_3)}}};
        CtrlState_dataBuf <= rndFuc_io_result;
      end else begin
        if(CtrlState_ongoing) begin
          CtrlState_enginRdy <= 1'b0;
          CtrlState_nextrndKey <= {_zz_CtrlState_nextrndKey_313,{_zz_CtrlState_nextrndKey_314,{_zz_CtrlState_nextrndKey_315,(_zz_CtrlState_nextrndKey_316 ^ _zz_CtrlState_nextrndKey_315)}}};
          CtrlState_dataBuf <= rndFuc_io_result;
          if(when_AES_CORE_l78) begin
            CtrlState_rndCnt <= (CtrlState_rndCnt + 4'b0001);
            CtrlState_ongoing <= 1'b1;
          end else begin
            CtrlState_rndCnt <= 4'b0000;
            CtrlState_ongoing <= 1'b0;
          end
        end else begin
          CtrlState_enginRdy <= 1'b1;
        end
      end
      CtrlState_lastRound_regNext <= CtrlState_lastRound;
    end
  end


endmodule
