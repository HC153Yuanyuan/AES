// Generator : SpinalHDL v1.7.0    git head : eca519e78d4e6022e34911ec300a432ed9db8220
// Component : MyroundFunction

`timescale 1ns/1ps 
module MyroundFunction (
  input      [127:0]  io_roundData,
  input               io_needMix,
  output     [127:0]  io_result
);

  wire       [31:0]   _zz_io_result;
  wire       [31:0]   _zz_io_result_1;
  wire       [31:0]   _zz_io_result_2;
  wire       [31:0]   _zz_io_result_3;
  reg        [31:0]   _zz_io_result_4;
  reg        [31:0]   _zz_io_result_5;
  reg        [31:0]   _zz_io_result_6;
  reg        [31:0]   _zz_io_result_7;
  reg        [31:0]   _zz_io_result_8;
  wire       [7:0]    _zz_io_result_9;
  reg        [7:0]    _zz_io_result_10;
  wire       [7:0]    _zz_io_result_11;
  reg        [7:0]    _zz_io_result_12;
  wire       [7:0]    _zz_io_result_13;
  reg        [7:0]    _zz_io_result_14;
  wire       [3:0]    _zz_io_result_15;
  wire       [3:0]    _zz_io_result_16;
  wire       [3:0]    _zz_io_result_17;
  reg        [3:0]    _zz_io_result_18;
  reg        [3:0]    _zz_io_result_19;
  wire       [1:0]    _zz_io_result_20;
  wire       [1:0]    _zz_io_result_21;
  wire       [1:0]    _zz_io_result_22;
  wire       [1:0]    _zz_io_result_23;
  wire       [1:0]    _zz_io_result_24;
  wire       [1:0]    _zz_io_result_25;
  wire       [1:0]    _zz_io_result_26;
  wire                _zz_io_result_27;
  reg        [1:0]    _zz_io_result_28;
  wire       [1:0]    _zz_io_result_29;
  reg        [1:0]    _zz_io_result_30;
  wire                _zz_io_result_31;
  reg        [1:0]    _zz_io_result_32;
  wire                _zz_io_result_33;
  reg        [1:0]    _zz_io_result_34;
  wire       [3:0]    _zz_io_result_35;
  wire       [3:0]    _zz_io_result_36;
  reg        [3:0]    _zz_io_result_37;
  wire       [1:0]    _zz_io_result_38;
  wire       [1:0]    _zz_io_result_39;
  wire       [1:0]    _zz_io_result_40;
  reg        [1:0]    _zz_io_result_41;
  wire                _zz_io_result_42;
  reg        [1:0]    _zz_io_result_43;
  wire       [1:0]    _zz_io_result_44;
  wire       [1:0]    _zz_io_result_45;
  reg        [1:0]    _zz_io_result_46;
  wire                _zz_io_result_47;
  reg        [1:0]    _zz_io_result_48;
  wire                _zz_io_result_49;
  reg        [1:0]    _zz_io_result_50;
  reg        [3:0]    _zz_io_result_51;
  wire       [1:0]    _zz_io_result_52;
  wire       [1:0]    _zz_io_result_53;
  wire       [1:0]    _zz_io_result_54;
  wire       [1:0]    _zz_io_result_55;
  wire       [1:0]    _zz_io_result_56;
  wire       [1:0]    _zz_io_result_57;
  wire       [1:0]    _zz_io_result_58;
  wire                _zz_io_result_59;
  reg        [1:0]    _zz_io_result_60;
  wire       [1:0]    _zz_io_result_61;
  reg        [1:0]    _zz_io_result_62;
  wire                _zz_io_result_63;
  reg        [1:0]    _zz_io_result_64;
  wire                _zz_io_result_65;
  reg        [1:0]    _zz_io_result_66;
  reg        [3:0]    _zz_io_result_67;
  wire       [1:0]    _zz_io_result_68;
  wire       [1:0]    _zz_io_result_69;
  wire       [1:0]    _zz_io_result_70;
  wire       [1:0]    _zz_io_result_71;
  wire       [1:0]    _zz_io_result_72;
  wire       [1:0]    _zz_io_result_73;
  wire       [1:0]    _zz_io_result_74;
  wire                _zz_io_result_75;
  reg        [1:0]    _zz_io_result_76;
  wire       [1:0]    _zz_io_result_77;
  reg        [1:0]    _zz_io_result_78;
  wire                _zz_io_result_79;
  reg        [1:0]    _zz_io_result_80;
  wire                _zz_io_result_81;
  reg        [1:0]    _zz_io_result_82;
  wire       [7:0]    _zz_io_result_83;
  reg        [7:0]    _zz_io_result_84;
  wire       [7:0]    _zz_io_result_85;
  reg        [7:0]    _zz_io_result_86;
  wire       [7:0]    _zz_io_result_87;
  reg        [7:0]    _zz_io_result_88;
  wire       [7:0]    _zz_io_result_89;
  reg        [7:0]    _zz_io_result_90;
  wire       [3:0]    _zz_io_result_91;
  wire       [3:0]    _zz_io_result_92;
  wire       [3:0]    _zz_io_result_93;
  reg        [3:0]    _zz_io_result_94;
  reg        [3:0]    _zz_io_result_95;
  wire       [1:0]    _zz_io_result_96;
  wire       [1:0]    _zz_io_result_97;
  wire       [1:0]    _zz_io_result_98;
  wire       [1:0]    _zz_io_result_99;
  wire       [1:0]    _zz_io_result_100;
  wire       [1:0]    _zz_io_result_101;
  wire       [1:0]    _zz_io_result_102;
  wire                _zz_io_result_103;
  reg        [1:0]    _zz_io_result_104;
  wire       [1:0]    _zz_io_result_105;
  reg        [1:0]    _zz_io_result_106;
  wire                _zz_io_result_107;
  reg        [1:0]    _zz_io_result_108;
  wire                _zz_io_result_109;
  reg        [1:0]    _zz_io_result_110;
  wire       [3:0]    _zz_io_result_111;
  wire       [3:0]    _zz_io_result_112;
  reg        [3:0]    _zz_io_result_113;
  wire       [1:0]    _zz_io_result_114;
  wire       [1:0]    _zz_io_result_115;
  wire       [1:0]    _zz_io_result_116;
  reg        [1:0]    _zz_io_result_117;
  wire                _zz_io_result_118;
  reg        [1:0]    _zz_io_result_119;
  wire       [1:0]    _zz_io_result_120;
  wire       [1:0]    _zz_io_result_121;
  reg        [1:0]    _zz_io_result_122;
  wire                _zz_io_result_123;
  reg        [1:0]    _zz_io_result_124;
  wire                _zz_io_result_125;
  reg        [1:0]    _zz_io_result_126;
  reg        [3:0]    _zz_io_result_127;
  wire       [1:0]    _zz_io_result_128;
  wire       [1:0]    _zz_io_result_129;
  wire       [1:0]    _zz_io_result_130;
  wire       [1:0]    _zz_io_result_131;
  wire       [1:0]    _zz_io_result_132;
  wire       [1:0]    _zz_io_result_133;
  wire       [1:0]    _zz_io_result_134;
  wire                _zz_io_result_135;
  reg        [1:0]    _zz_io_result_136;
  wire       [1:0]    _zz_io_result_137;
  reg        [1:0]    _zz_io_result_138;
  wire                _zz_io_result_139;
  reg        [1:0]    _zz_io_result_140;
  wire                _zz_io_result_141;
  reg        [1:0]    _zz_io_result_142;
  reg        [3:0]    _zz_io_result_143;
  wire       [1:0]    _zz_io_result_144;
  wire       [1:0]    _zz_io_result_145;
  wire       [1:0]    _zz_io_result_146;
  wire       [1:0]    _zz_io_result_147;
  wire       [1:0]    _zz_io_result_148;
  wire       [1:0]    _zz_io_result_149;
  wire       [1:0]    _zz_io_result_150;
  wire                _zz_io_result_151;
  reg        [1:0]    _zz_io_result_152;
  wire       [1:0]    _zz_io_result_153;
  reg        [1:0]    _zz_io_result_154;
  wire                _zz_io_result_155;
  reg        [1:0]    _zz_io_result_156;
  wire                _zz_io_result_157;
  reg        [1:0]    _zz_io_result_158;
  wire       [7:0]    _zz_io_result_159;
  reg        [7:0]    _zz_io_result_160;
  wire       [7:0]    _zz_io_result_161;
  reg        [7:0]    _zz_io_result_162;
  wire       [7:0]    _zz_io_result_163;
  reg        [7:0]    _zz_io_result_164;
  wire       [7:0]    _zz_io_result_165;
  reg        [7:0]    _zz_io_result_166;
  wire       [3:0]    _zz_io_result_167;
  wire       [3:0]    _zz_io_result_168;
  wire       [3:0]    _zz_io_result_169;
  reg        [3:0]    _zz_io_result_170;
  reg        [3:0]    _zz_io_result_171;
  wire       [1:0]    _zz_io_result_172;
  wire       [1:0]    _zz_io_result_173;
  wire       [1:0]    _zz_io_result_174;
  wire       [1:0]    _zz_io_result_175;
  wire       [1:0]    _zz_io_result_176;
  wire       [1:0]    _zz_io_result_177;
  wire       [1:0]    _zz_io_result_178;
  wire                _zz_io_result_179;
  reg        [1:0]    _zz_io_result_180;
  wire       [1:0]    _zz_io_result_181;
  reg        [1:0]    _zz_io_result_182;
  wire                _zz_io_result_183;
  reg        [1:0]    _zz_io_result_184;
  wire                _zz_io_result_185;
  reg        [1:0]    _zz_io_result_186;
  wire       [3:0]    _zz_io_result_187;
  wire       [3:0]    _zz_io_result_188;
  reg        [3:0]    _zz_io_result_189;
  wire       [1:0]    _zz_io_result_190;
  wire       [1:0]    _zz_io_result_191;
  wire       [1:0]    _zz_io_result_192;
  reg        [1:0]    _zz_io_result_193;
  wire                _zz_io_result_194;
  reg        [1:0]    _zz_io_result_195;
  wire       [1:0]    _zz_io_result_196;
  wire       [1:0]    _zz_io_result_197;
  reg        [1:0]    _zz_io_result_198;
  wire                _zz_io_result_199;
  reg        [1:0]    _zz_io_result_200;
  wire                _zz_io_result_201;
  reg        [1:0]    _zz_io_result_202;
  reg        [3:0]    _zz_io_result_203;
  wire       [1:0]    _zz_io_result_204;
  wire       [1:0]    _zz_io_result_205;
  wire       [1:0]    _zz_io_result_206;
  wire       [1:0]    _zz_io_result_207;
  wire       [1:0]    _zz_io_result_208;
  wire       [1:0]    _zz_io_result_209;
  wire       [1:0]    _zz_io_result_210;
  wire                _zz_io_result_211;
  reg        [1:0]    _zz_io_result_212;
  wire       [1:0]    _zz_io_result_213;
  reg        [1:0]    _zz_io_result_214;
  wire                _zz_io_result_215;
  reg        [1:0]    _zz_io_result_216;
  wire                _zz_io_result_217;
  reg        [1:0]    _zz_io_result_218;
  reg        [3:0]    _zz_io_result_219;
  wire       [1:0]    _zz_io_result_220;
  wire       [1:0]    _zz_io_result_221;
  wire       [1:0]    _zz_io_result_222;
  wire       [1:0]    _zz_io_result_223;
  wire       [1:0]    _zz_io_result_224;
  wire       [1:0]    _zz_io_result_225;
  wire       [1:0]    _zz_io_result_226;
  wire                _zz_io_result_227;
  reg        [1:0]    _zz_io_result_228;
  wire       [1:0]    _zz_io_result_229;
  reg        [1:0]    _zz_io_result_230;
  wire                _zz_io_result_231;
  reg        [1:0]    _zz_io_result_232;
  wire                _zz_io_result_233;
  reg        [1:0]    _zz_io_result_234;
  wire       [7:0]    _zz_io_result_235;
  reg        [7:0]    _zz_io_result_236;
  wire       [7:0]    _zz_io_result_237;
  reg        [7:0]    _zz_io_result_238;
  wire       [7:0]    _zz_io_result_239;
  reg        [7:0]    _zz_io_result_240;
  wire       [7:0]    _zz_io_result_241;
  reg        [7:0]    _zz_io_result_242;
  wire       [3:0]    _zz_io_result_243;
  wire       [3:0]    _zz_io_result_244;
  wire       [3:0]    _zz_io_result_245;
  reg        [3:0]    _zz_io_result_246;
  reg        [3:0]    _zz_io_result_247;
  wire       [1:0]    _zz_io_result_248;
  wire       [1:0]    _zz_io_result_249;
  wire       [1:0]    _zz_io_result_250;
  wire       [1:0]    _zz_io_result_251;
  wire       [1:0]    _zz_io_result_252;
  wire       [1:0]    _zz_io_result_253;
  wire       [1:0]    _zz_io_result_254;
  wire                _zz_io_result_255;
  reg        [1:0]    _zz_io_result_256;
  wire       [1:0]    _zz_io_result_257;
  reg        [1:0]    _zz_io_result_258;
  wire                _zz_io_result_259;
  reg        [1:0]    _zz_io_result_260;
  wire                _zz_io_result_261;
  reg        [1:0]    _zz_io_result_262;
  wire       [3:0]    _zz_io_result_263;
  wire       [3:0]    _zz_io_result_264;
  reg        [3:0]    _zz_io_result_265;
  wire       [1:0]    _zz_io_result_266;
  wire       [1:0]    _zz_io_result_267;
  wire       [1:0]    _zz_io_result_268;
  reg        [1:0]    _zz_io_result_269;
  wire                _zz_io_result_270;
  reg        [1:0]    _zz_io_result_271;
  wire       [1:0]    _zz_io_result_272;
  wire       [1:0]    _zz_io_result_273;
  reg        [1:0]    _zz_io_result_274;
  wire                _zz_io_result_275;
  reg        [1:0]    _zz_io_result_276;
  wire                _zz_io_result_277;
  reg        [1:0]    _zz_io_result_278;
  reg        [3:0]    _zz_io_result_279;
  wire       [1:0]    _zz_io_result_280;
  wire       [1:0]    _zz_io_result_281;
  wire       [1:0]    _zz_io_result_282;
  wire       [1:0]    _zz_io_result_283;
  wire       [1:0]    _zz_io_result_284;
  wire       [1:0]    _zz_io_result_285;
  wire       [1:0]    _zz_io_result_286;
  wire                _zz_io_result_287;
  reg        [1:0]    _zz_io_result_288;
  wire       [1:0]    _zz_io_result_289;
  reg        [1:0]    _zz_io_result_290;
  wire                _zz_io_result_291;
  reg        [1:0]    _zz_io_result_292;
  wire                _zz_io_result_293;
  reg        [1:0]    _zz_io_result_294;
  reg        [3:0]    _zz_io_result_295;
  wire       [1:0]    _zz_io_result_296;
  wire       [1:0]    _zz_io_result_297;
  wire       [1:0]    _zz_io_result_298;
  wire       [1:0]    _zz_io_result_299;
  wire       [1:0]    _zz_io_result_300;
  wire       [1:0]    _zz_io_result_301;
  wire       [1:0]    _zz_io_result_302;
  wire                _zz_io_result_303;
  reg        [1:0]    _zz_io_result_304;
  wire       [1:0]    _zz_io_result_305;
  reg        [1:0]    _zz_io_result_306;
  wire                _zz_io_result_307;
  reg        [1:0]    _zz_io_result_308;
  wire                _zz_io_result_309;
  reg        [1:0]    _zz_io_result_310;
  wire       [7:0]    _zz_io_result_311;
  reg        [7:0]    _zz_io_result_312;
  reg        [31:0]   _zz_io_result_313;
  wire       [7:0]    _zz_io_result_314;
  reg        [7:0]    _zz_io_result_315;
  wire       [7:0]    _zz_io_result_316;
  reg        [7:0]    _zz_io_result_317;
  wire       [7:0]    _zz_io_result_318;
  reg        [7:0]    _zz_io_result_319;
  wire       [3:0]    _zz_io_result_320;
  wire       [3:0]    _zz_io_result_321;
  wire       [3:0]    _zz_io_result_322;
  reg        [3:0]    _zz_io_result_323;
  reg        [3:0]    _zz_io_result_324;
  wire       [1:0]    _zz_io_result_325;
  wire       [1:0]    _zz_io_result_326;
  wire       [1:0]    _zz_io_result_327;
  wire       [1:0]    _zz_io_result_328;
  wire       [1:0]    _zz_io_result_329;
  wire       [1:0]    _zz_io_result_330;
  wire       [1:0]    _zz_io_result_331;
  wire                _zz_io_result_332;
  reg        [1:0]    _zz_io_result_333;
  wire       [1:0]    _zz_io_result_334;
  reg        [1:0]    _zz_io_result_335;
  wire                _zz_io_result_336;
  reg        [1:0]    _zz_io_result_337;
  wire                _zz_io_result_338;
  reg        [1:0]    _zz_io_result_339;
  wire       [3:0]    _zz_io_result_340;
  wire       [3:0]    _zz_io_result_341;
  reg        [3:0]    _zz_io_result_342;
  wire       [1:0]    _zz_io_result_343;
  wire       [1:0]    _zz_io_result_344;
  wire       [1:0]    _zz_io_result_345;
  reg        [1:0]    _zz_io_result_346;
  wire                _zz_io_result_347;
  reg        [1:0]    _zz_io_result_348;
  wire       [1:0]    _zz_io_result_349;
  wire       [1:0]    _zz_io_result_350;
  reg        [1:0]    _zz_io_result_351;
  wire                _zz_io_result_352;
  reg        [1:0]    _zz_io_result_353;
  wire                _zz_io_result_354;
  reg        [1:0]    _zz_io_result_355;
  reg        [3:0]    _zz_io_result_356;
  wire       [1:0]    _zz_io_result_357;
  wire       [1:0]    _zz_io_result_358;
  wire       [1:0]    _zz_io_result_359;
  wire       [1:0]    _zz_io_result_360;
  wire       [1:0]    _zz_io_result_361;
  wire       [1:0]    _zz_io_result_362;
  wire       [1:0]    _zz_io_result_363;
  wire                _zz_io_result_364;
  reg        [1:0]    _zz_io_result_365;
  wire       [1:0]    _zz_io_result_366;
  reg        [1:0]    _zz_io_result_367;
  wire                _zz_io_result_368;
  reg        [1:0]    _zz_io_result_369;
  wire                _zz_io_result_370;
  reg        [1:0]    _zz_io_result_371;
  reg        [3:0]    _zz_io_result_372;
  wire       [1:0]    _zz_io_result_373;
  wire       [1:0]    _zz_io_result_374;
  wire       [1:0]    _zz_io_result_375;
  wire       [1:0]    _zz_io_result_376;
  wire       [1:0]    _zz_io_result_377;
  wire       [1:0]    _zz_io_result_378;
  wire       [1:0]    _zz_io_result_379;
  wire                _zz_io_result_380;
  reg        [1:0]    _zz_io_result_381;
  wire       [1:0]    _zz_io_result_382;
  reg        [1:0]    _zz_io_result_383;
  wire                _zz_io_result_384;
  reg        [1:0]    _zz_io_result_385;
  wire                _zz_io_result_386;
  reg        [1:0]    _zz_io_result_387;
  wire       [7:0]    _zz_io_result_388;
  reg        [7:0]    _zz_io_result_389;
  wire       [7:0]    _zz_io_result_390;
  reg        [7:0]    _zz_io_result_391;
  wire       [7:0]    _zz_io_result_392;
  reg        [7:0]    _zz_io_result_393;
  wire       [7:0]    _zz_io_result_394;
  reg        [7:0]    _zz_io_result_395;
  wire       [3:0]    _zz_io_result_396;
  wire       [3:0]    _zz_io_result_397;
  wire       [3:0]    _zz_io_result_398;
  reg        [3:0]    _zz_io_result_399;
  reg        [3:0]    _zz_io_result_400;
  wire       [1:0]    _zz_io_result_401;
  wire       [1:0]    _zz_io_result_402;
  wire       [1:0]    _zz_io_result_403;
  wire       [1:0]    _zz_io_result_404;
  wire       [1:0]    _zz_io_result_405;
  wire       [1:0]    _zz_io_result_406;
  wire       [1:0]    _zz_io_result_407;
  wire                _zz_io_result_408;
  reg        [1:0]    _zz_io_result_409;
  wire       [1:0]    _zz_io_result_410;
  reg        [1:0]    _zz_io_result_411;
  wire                _zz_io_result_412;
  reg        [1:0]    _zz_io_result_413;
  wire                _zz_io_result_414;
  reg        [1:0]    _zz_io_result_415;
  wire       [3:0]    _zz_io_result_416;
  wire       [3:0]    _zz_io_result_417;
  reg        [3:0]    _zz_io_result_418;
  wire       [1:0]    _zz_io_result_419;
  wire       [1:0]    _zz_io_result_420;
  wire       [1:0]    _zz_io_result_421;
  reg        [1:0]    _zz_io_result_422;
  wire                _zz_io_result_423;
  reg        [1:0]    _zz_io_result_424;
  wire       [1:0]    _zz_io_result_425;
  wire       [1:0]    _zz_io_result_426;
  reg        [1:0]    _zz_io_result_427;
  wire                _zz_io_result_428;
  reg        [1:0]    _zz_io_result_429;
  wire                _zz_io_result_430;
  reg        [1:0]    _zz_io_result_431;
  reg        [3:0]    _zz_io_result_432;
  wire       [1:0]    _zz_io_result_433;
  wire       [1:0]    _zz_io_result_434;
  wire       [1:0]    _zz_io_result_435;
  wire       [1:0]    _zz_io_result_436;
  wire       [1:0]    _zz_io_result_437;
  wire       [1:0]    _zz_io_result_438;
  wire       [1:0]    _zz_io_result_439;
  wire                _zz_io_result_440;
  reg        [1:0]    _zz_io_result_441;
  wire       [1:0]    _zz_io_result_442;
  reg        [1:0]    _zz_io_result_443;
  wire                _zz_io_result_444;
  reg        [1:0]    _zz_io_result_445;
  wire                _zz_io_result_446;
  reg        [1:0]    _zz_io_result_447;
  reg        [3:0]    _zz_io_result_448;
  wire       [1:0]    _zz_io_result_449;
  wire       [1:0]    _zz_io_result_450;
  wire       [1:0]    _zz_io_result_451;
  wire       [1:0]    _zz_io_result_452;
  wire       [1:0]    _zz_io_result_453;
  wire       [1:0]    _zz_io_result_454;
  wire       [1:0]    _zz_io_result_455;
  wire                _zz_io_result_456;
  reg        [1:0]    _zz_io_result_457;
  wire       [1:0]    _zz_io_result_458;
  reg        [1:0]    _zz_io_result_459;
  wire                _zz_io_result_460;
  reg        [1:0]    _zz_io_result_461;
  wire                _zz_io_result_462;
  reg        [1:0]    _zz_io_result_463;
  wire       [7:0]    _zz_io_result_464;
  reg        [7:0]    _zz_io_result_465;
  wire       [7:0]    _zz_io_result_466;
  reg        [7:0]    _zz_io_result_467;
  wire       [7:0]    _zz_io_result_468;
  reg        [7:0]    _zz_io_result_469;
  wire       [7:0]    _zz_io_result_470;
  reg        [7:0]    _zz_io_result_471;
  wire       [3:0]    _zz_io_result_472;
  wire       [3:0]    _zz_io_result_473;
  wire       [3:0]    _zz_io_result_474;
  reg        [3:0]    _zz_io_result_475;
  reg        [3:0]    _zz_io_result_476;
  wire       [1:0]    _zz_io_result_477;
  wire       [1:0]    _zz_io_result_478;
  wire       [1:0]    _zz_io_result_479;
  wire       [1:0]    _zz_io_result_480;
  wire       [1:0]    _zz_io_result_481;
  wire       [1:0]    _zz_io_result_482;
  wire       [1:0]    _zz_io_result_483;
  wire                _zz_io_result_484;
  reg        [1:0]    _zz_io_result_485;
  wire       [1:0]    _zz_io_result_486;
  reg        [1:0]    _zz_io_result_487;
  wire                _zz_io_result_488;
  reg        [1:0]    _zz_io_result_489;
  wire                _zz_io_result_490;
  reg        [1:0]    _zz_io_result_491;
  wire       [3:0]    _zz_io_result_492;
  wire       [3:0]    _zz_io_result_493;
  reg        [3:0]    _zz_io_result_494;
  wire       [1:0]    _zz_io_result_495;
  wire       [1:0]    _zz_io_result_496;
  wire       [1:0]    _zz_io_result_497;
  reg        [1:0]    _zz_io_result_498;
  wire                _zz_io_result_499;
  reg        [1:0]    _zz_io_result_500;
  wire       [1:0]    _zz_io_result_501;
  wire       [1:0]    _zz_io_result_502;
  reg        [1:0]    _zz_io_result_503;
  wire                _zz_io_result_504;
  reg        [1:0]    _zz_io_result_505;
  wire                _zz_io_result_506;
  reg        [1:0]    _zz_io_result_507;
  reg        [3:0]    _zz_io_result_508;
  wire       [1:0]    _zz_io_result_509;
  wire       [1:0]    _zz_io_result_510;
  wire       [1:0]    _zz_io_result_511;
  wire       [1:0]    _zz_io_result_512;
  wire       [1:0]    _zz_io_result_513;
  wire       [1:0]    _zz_io_result_514;
  wire       [1:0]    _zz_io_result_515;
  wire                _zz_io_result_516;
  reg        [1:0]    _zz_io_result_517;
  wire       [1:0]    _zz_io_result_518;
  reg        [1:0]    _zz_io_result_519;
  wire                _zz_io_result_520;
  reg        [1:0]    _zz_io_result_521;
  wire                _zz_io_result_522;
  reg        [1:0]    _zz_io_result_523;
  reg        [3:0]    _zz_io_result_524;
  wire       [1:0]    _zz_io_result_525;
  wire       [1:0]    _zz_io_result_526;
  wire       [1:0]    _zz_io_result_527;
  wire       [1:0]    _zz_io_result_528;
  wire       [1:0]    _zz_io_result_529;
  wire       [1:0]    _zz_io_result_530;
  wire       [1:0]    _zz_io_result_531;
  wire                _zz_io_result_532;
  reg        [1:0]    _zz_io_result_533;
  wire       [1:0]    _zz_io_result_534;
  reg        [1:0]    _zz_io_result_535;
  wire                _zz_io_result_536;
  reg        [1:0]    _zz_io_result_537;
  wire                _zz_io_result_538;
  reg        [1:0]    _zz_io_result_539;
  wire       [7:0]    _zz_io_result_540;
  reg        [7:0]    _zz_io_result_541;
  wire       [7:0]    _zz_io_result_542;
  reg        [7:0]    _zz_io_result_543;
  wire       [7:0]    _zz_io_result_544;
  reg        [7:0]    _zz_io_result_545;
  wire       [7:0]    _zz_io_result_546;
  reg        [7:0]    _zz_io_result_547;
  wire       [3:0]    _zz_io_result_548;
  wire       [3:0]    _zz_io_result_549;
  wire       [3:0]    _zz_io_result_550;
  reg        [3:0]    _zz_io_result_551;
  reg        [3:0]    _zz_io_result_552;
  wire       [1:0]    _zz_io_result_553;
  wire       [1:0]    _zz_io_result_554;
  wire       [1:0]    _zz_io_result_555;
  wire       [1:0]    _zz_io_result_556;
  wire       [1:0]    _zz_io_result_557;
  wire       [1:0]    _zz_io_result_558;
  wire       [1:0]    _zz_io_result_559;
  wire                _zz_io_result_560;
  reg        [1:0]    _zz_io_result_561;
  wire       [1:0]    _zz_io_result_562;
  reg        [1:0]    _zz_io_result_563;
  wire                _zz_io_result_564;
  reg        [1:0]    _zz_io_result_565;
  wire                _zz_io_result_566;
  reg        [1:0]    _zz_io_result_567;
  wire       [3:0]    _zz_io_result_568;
  wire       [3:0]    _zz_io_result_569;
  reg        [3:0]    _zz_io_result_570;
  wire       [1:0]    _zz_io_result_571;
  wire       [1:0]    _zz_io_result_572;
  wire       [1:0]    _zz_io_result_573;
  reg        [1:0]    _zz_io_result_574;
  wire                _zz_io_result_575;
  reg        [1:0]    _zz_io_result_576;
  wire       [1:0]    _zz_io_result_577;
  wire       [1:0]    _zz_io_result_578;
  reg        [1:0]    _zz_io_result_579;
  wire                _zz_io_result_580;
  reg        [1:0]    _zz_io_result_581;
  wire                _zz_io_result_582;
  reg        [1:0]    _zz_io_result_583;
  reg        [3:0]    _zz_io_result_584;
  wire       [1:0]    _zz_io_result_585;
  wire       [1:0]    _zz_io_result_586;
  wire       [1:0]    _zz_io_result_587;
  wire       [1:0]    _zz_io_result_588;
  wire       [1:0]    _zz_io_result_589;
  wire       [1:0]    _zz_io_result_590;
  wire       [1:0]    _zz_io_result_591;
  wire                _zz_io_result_592;
  reg        [1:0]    _zz_io_result_593;
  wire       [1:0]    _zz_io_result_594;
  reg        [1:0]    _zz_io_result_595;
  wire                _zz_io_result_596;
  reg        [1:0]    _zz_io_result_597;
  wire                _zz_io_result_598;
  reg        [1:0]    _zz_io_result_599;
  reg        [3:0]    _zz_io_result_600;
  wire       [1:0]    _zz_io_result_601;
  wire       [1:0]    _zz_io_result_602;
  wire       [1:0]    _zz_io_result_603;
  wire       [1:0]    _zz_io_result_604;
  wire       [1:0]    _zz_io_result_605;
  wire       [1:0]    _zz_io_result_606;
  wire       [1:0]    _zz_io_result_607;
  wire                _zz_io_result_608;
  reg        [1:0]    _zz_io_result_609;
  wire       [1:0]    _zz_io_result_610;
  reg        [1:0]    _zz_io_result_611;
  wire                _zz_io_result_612;
  reg        [1:0]    _zz_io_result_613;
  wire                _zz_io_result_614;
  reg        [1:0]    _zz_io_result_615;
  wire       [7:0]    _zz_io_result_616;
  reg        [7:0]    _zz_io_result_617;
  reg        [31:0]   _zz_io_result_618;
  wire       [7:0]    _zz_io_result_619;
  reg        [7:0]    _zz_io_result_620;
  wire       [7:0]    _zz_io_result_621;
  reg        [7:0]    _zz_io_result_622;
  wire       [7:0]    _zz_io_result_623;
  reg        [7:0]    _zz_io_result_624;
  wire       [3:0]    _zz_io_result_625;
  wire       [3:0]    _zz_io_result_626;
  wire       [3:0]    _zz_io_result_627;
  reg        [3:0]    _zz_io_result_628;
  reg        [3:0]    _zz_io_result_629;
  wire       [1:0]    _zz_io_result_630;
  wire       [1:0]    _zz_io_result_631;
  wire       [1:0]    _zz_io_result_632;
  wire       [1:0]    _zz_io_result_633;
  wire       [1:0]    _zz_io_result_634;
  wire       [1:0]    _zz_io_result_635;
  wire       [1:0]    _zz_io_result_636;
  wire                _zz_io_result_637;
  reg        [1:0]    _zz_io_result_638;
  wire       [1:0]    _zz_io_result_639;
  reg        [1:0]    _zz_io_result_640;
  wire                _zz_io_result_641;
  reg        [1:0]    _zz_io_result_642;
  wire                _zz_io_result_643;
  reg        [1:0]    _zz_io_result_644;
  wire       [3:0]    _zz_io_result_645;
  wire       [3:0]    _zz_io_result_646;
  reg        [3:0]    _zz_io_result_647;
  wire       [1:0]    _zz_io_result_648;
  wire       [1:0]    _zz_io_result_649;
  wire       [1:0]    _zz_io_result_650;
  reg        [1:0]    _zz_io_result_651;
  wire                _zz_io_result_652;
  reg        [1:0]    _zz_io_result_653;
  wire       [1:0]    _zz_io_result_654;
  wire       [1:0]    _zz_io_result_655;
  reg        [1:0]    _zz_io_result_656;
  wire                _zz_io_result_657;
  reg        [1:0]    _zz_io_result_658;
  wire                _zz_io_result_659;
  reg        [1:0]    _zz_io_result_660;
  reg        [3:0]    _zz_io_result_661;
  wire       [1:0]    _zz_io_result_662;
  wire       [1:0]    _zz_io_result_663;
  wire       [1:0]    _zz_io_result_664;
  wire       [1:0]    _zz_io_result_665;
  wire       [1:0]    _zz_io_result_666;
  wire       [1:0]    _zz_io_result_667;
  wire       [1:0]    _zz_io_result_668;
  wire                _zz_io_result_669;
  reg        [1:0]    _zz_io_result_670;
  wire       [1:0]    _zz_io_result_671;
  reg        [1:0]    _zz_io_result_672;
  wire                _zz_io_result_673;
  reg        [1:0]    _zz_io_result_674;
  wire                _zz_io_result_675;
  reg        [1:0]    _zz_io_result_676;
  reg        [3:0]    _zz_io_result_677;
  wire       [1:0]    _zz_io_result_678;
  wire       [1:0]    _zz_io_result_679;
  wire       [1:0]    _zz_io_result_680;
  wire       [1:0]    _zz_io_result_681;
  wire       [1:0]    _zz_io_result_682;
  wire       [1:0]    _zz_io_result_683;
  wire       [1:0]    _zz_io_result_684;
  wire                _zz_io_result_685;
  reg        [1:0]    _zz_io_result_686;
  wire       [1:0]    _zz_io_result_687;
  reg        [1:0]    _zz_io_result_688;
  wire                _zz_io_result_689;
  reg        [1:0]    _zz_io_result_690;
  wire                _zz_io_result_691;
  reg        [1:0]    _zz_io_result_692;
  wire       [7:0]    _zz_io_result_693;
  reg        [7:0]    _zz_io_result_694;
  wire       [7:0]    _zz_io_result_695;
  reg        [7:0]    _zz_io_result_696;
  wire       [7:0]    _zz_io_result_697;
  reg        [7:0]    _zz_io_result_698;
  wire       [7:0]    _zz_io_result_699;
  reg        [7:0]    _zz_io_result_700;
  wire       [3:0]    _zz_io_result_701;
  wire       [3:0]    _zz_io_result_702;
  wire       [3:0]    _zz_io_result_703;
  reg        [3:0]    _zz_io_result_704;
  reg        [3:0]    _zz_io_result_705;
  wire       [1:0]    _zz_io_result_706;
  wire       [1:0]    _zz_io_result_707;
  wire       [1:0]    _zz_io_result_708;
  wire       [1:0]    _zz_io_result_709;
  wire       [1:0]    _zz_io_result_710;
  wire       [1:0]    _zz_io_result_711;
  wire       [1:0]    _zz_io_result_712;
  wire                _zz_io_result_713;
  reg        [1:0]    _zz_io_result_714;
  wire       [1:0]    _zz_io_result_715;
  reg        [1:0]    _zz_io_result_716;
  wire                _zz_io_result_717;
  reg        [1:0]    _zz_io_result_718;
  wire                _zz_io_result_719;
  reg        [1:0]    _zz_io_result_720;
  wire       [3:0]    _zz_io_result_721;
  wire       [3:0]    _zz_io_result_722;
  reg        [3:0]    _zz_io_result_723;
  wire       [1:0]    _zz_io_result_724;
  wire       [1:0]    _zz_io_result_725;
  wire       [1:0]    _zz_io_result_726;
  reg        [1:0]    _zz_io_result_727;
  wire                _zz_io_result_728;
  reg        [1:0]    _zz_io_result_729;
  wire       [1:0]    _zz_io_result_730;
  wire       [1:0]    _zz_io_result_731;
  reg        [1:0]    _zz_io_result_732;
  wire                _zz_io_result_733;
  reg        [1:0]    _zz_io_result_734;
  wire                _zz_io_result_735;
  reg        [1:0]    _zz_io_result_736;
  reg        [3:0]    _zz_io_result_737;
  wire       [1:0]    _zz_io_result_738;
  wire       [1:0]    _zz_io_result_739;
  wire       [1:0]    _zz_io_result_740;
  wire       [1:0]    _zz_io_result_741;
  wire       [1:0]    _zz_io_result_742;
  wire       [1:0]    _zz_io_result_743;
  wire       [1:0]    _zz_io_result_744;
  wire                _zz_io_result_745;
  reg        [1:0]    _zz_io_result_746;
  wire       [1:0]    _zz_io_result_747;
  reg        [1:0]    _zz_io_result_748;
  wire                _zz_io_result_749;
  reg        [1:0]    _zz_io_result_750;
  wire                _zz_io_result_751;
  reg        [1:0]    _zz_io_result_752;
  reg        [3:0]    _zz_io_result_753;
  wire       [1:0]    _zz_io_result_754;
  wire       [1:0]    _zz_io_result_755;
  wire       [1:0]    _zz_io_result_756;
  wire       [1:0]    _zz_io_result_757;
  wire       [1:0]    _zz_io_result_758;
  wire       [1:0]    _zz_io_result_759;
  wire       [1:0]    _zz_io_result_760;
  wire                _zz_io_result_761;
  reg        [1:0]    _zz_io_result_762;
  wire       [1:0]    _zz_io_result_763;
  reg        [1:0]    _zz_io_result_764;
  wire                _zz_io_result_765;
  reg        [1:0]    _zz_io_result_766;
  wire                _zz_io_result_767;
  reg        [1:0]    _zz_io_result_768;
  wire       [7:0]    _zz_io_result_769;
  reg        [7:0]    _zz_io_result_770;
  wire       [7:0]    _zz_io_result_771;
  reg        [7:0]    _zz_io_result_772;
  wire       [7:0]    _zz_io_result_773;
  reg        [7:0]    _zz_io_result_774;
  wire       [7:0]    _zz_io_result_775;
  reg        [7:0]    _zz_io_result_776;
  wire       [3:0]    _zz_io_result_777;
  wire       [3:0]    _zz_io_result_778;
  wire       [3:0]    _zz_io_result_779;
  reg        [3:0]    _zz_io_result_780;
  reg        [3:0]    _zz_io_result_781;
  wire       [1:0]    _zz_io_result_782;
  wire       [1:0]    _zz_io_result_783;
  wire       [1:0]    _zz_io_result_784;
  wire       [1:0]    _zz_io_result_785;
  wire       [1:0]    _zz_io_result_786;
  wire       [1:0]    _zz_io_result_787;
  wire       [1:0]    _zz_io_result_788;
  wire                _zz_io_result_789;
  reg        [1:0]    _zz_io_result_790;
  wire       [1:0]    _zz_io_result_791;
  reg        [1:0]    _zz_io_result_792;
  wire                _zz_io_result_793;
  reg        [1:0]    _zz_io_result_794;
  wire                _zz_io_result_795;
  reg        [1:0]    _zz_io_result_796;
  wire       [3:0]    _zz_io_result_797;
  wire       [3:0]    _zz_io_result_798;
  reg        [3:0]    _zz_io_result_799;
  wire       [1:0]    _zz_io_result_800;
  wire       [1:0]    _zz_io_result_801;
  wire       [1:0]    _zz_io_result_802;
  reg        [1:0]    _zz_io_result_803;
  wire                _zz_io_result_804;
  reg        [1:0]    _zz_io_result_805;
  wire       [1:0]    _zz_io_result_806;
  wire       [1:0]    _zz_io_result_807;
  reg        [1:0]    _zz_io_result_808;
  wire                _zz_io_result_809;
  reg        [1:0]    _zz_io_result_810;
  wire                _zz_io_result_811;
  reg        [1:0]    _zz_io_result_812;
  reg        [3:0]    _zz_io_result_813;
  wire       [1:0]    _zz_io_result_814;
  wire       [1:0]    _zz_io_result_815;
  wire       [1:0]    _zz_io_result_816;
  wire       [1:0]    _zz_io_result_817;
  wire       [1:0]    _zz_io_result_818;
  wire       [1:0]    _zz_io_result_819;
  wire       [1:0]    _zz_io_result_820;
  wire                _zz_io_result_821;
  reg        [1:0]    _zz_io_result_822;
  wire       [1:0]    _zz_io_result_823;
  reg        [1:0]    _zz_io_result_824;
  wire                _zz_io_result_825;
  reg        [1:0]    _zz_io_result_826;
  wire                _zz_io_result_827;
  reg        [1:0]    _zz_io_result_828;
  reg        [3:0]    _zz_io_result_829;
  wire       [1:0]    _zz_io_result_830;
  wire       [1:0]    _zz_io_result_831;
  wire       [1:0]    _zz_io_result_832;
  wire       [1:0]    _zz_io_result_833;
  wire       [1:0]    _zz_io_result_834;
  wire       [1:0]    _zz_io_result_835;
  wire       [1:0]    _zz_io_result_836;
  wire                _zz_io_result_837;
  reg        [1:0]    _zz_io_result_838;
  wire       [1:0]    _zz_io_result_839;
  reg        [1:0]    _zz_io_result_840;
  wire                _zz_io_result_841;
  reg        [1:0]    _zz_io_result_842;
  wire                _zz_io_result_843;
  reg        [1:0]    _zz_io_result_844;
  wire       [7:0]    _zz_io_result_845;
  reg        [7:0]    _zz_io_result_846;
  wire       [7:0]    _zz_io_result_847;
  reg        [7:0]    _zz_io_result_848;
  wire       [7:0]    _zz_io_result_849;
  reg        [7:0]    _zz_io_result_850;
  wire       [7:0]    _zz_io_result_851;
  reg        [7:0]    _zz_io_result_852;
  wire       [3:0]    _zz_io_result_853;
  wire       [3:0]    _zz_io_result_854;
  wire       [3:0]    _zz_io_result_855;
  reg        [3:0]    _zz_io_result_856;
  reg        [3:0]    _zz_io_result_857;
  wire       [1:0]    _zz_io_result_858;
  wire       [1:0]    _zz_io_result_859;
  wire       [1:0]    _zz_io_result_860;
  wire       [1:0]    _zz_io_result_861;
  wire       [1:0]    _zz_io_result_862;
  wire       [1:0]    _zz_io_result_863;
  wire       [1:0]    _zz_io_result_864;
  wire                _zz_io_result_865;
  reg        [1:0]    _zz_io_result_866;
  wire       [1:0]    _zz_io_result_867;
  reg        [1:0]    _zz_io_result_868;
  wire                _zz_io_result_869;
  reg        [1:0]    _zz_io_result_870;
  wire                _zz_io_result_871;
  reg        [1:0]    _zz_io_result_872;
  wire       [3:0]    _zz_io_result_873;
  wire       [3:0]    _zz_io_result_874;
  reg        [3:0]    _zz_io_result_875;
  wire       [1:0]    _zz_io_result_876;
  wire       [1:0]    _zz_io_result_877;
  wire       [1:0]    _zz_io_result_878;
  reg        [1:0]    _zz_io_result_879;
  wire                _zz_io_result_880;
  reg        [1:0]    _zz_io_result_881;
  wire       [1:0]    _zz_io_result_882;
  wire       [1:0]    _zz_io_result_883;
  reg        [1:0]    _zz_io_result_884;
  wire                _zz_io_result_885;
  reg        [1:0]    _zz_io_result_886;
  wire                _zz_io_result_887;
  reg        [1:0]    _zz_io_result_888;
  reg        [3:0]    _zz_io_result_889;
  wire       [1:0]    _zz_io_result_890;
  wire       [1:0]    _zz_io_result_891;
  wire       [1:0]    _zz_io_result_892;
  wire       [1:0]    _zz_io_result_893;
  wire       [1:0]    _zz_io_result_894;
  wire       [1:0]    _zz_io_result_895;
  wire       [1:0]    _zz_io_result_896;
  wire                _zz_io_result_897;
  reg        [1:0]    _zz_io_result_898;
  wire       [1:0]    _zz_io_result_899;
  reg        [1:0]    _zz_io_result_900;
  wire                _zz_io_result_901;
  reg        [1:0]    _zz_io_result_902;
  wire                _zz_io_result_903;
  reg        [1:0]    _zz_io_result_904;
  reg        [3:0]    _zz_io_result_905;
  wire       [1:0]    _zz_io_result_906;
  wire       [1:0]    _zz_io_result_907;
  wire       [1:0]    _zz_io_result_908;
  wire       [1:0]    _zz_io_result_909;
  wire       [1:0]    _zz_io_result_910;
  wire       [1:0]    _zz_io_result_911;
  wire       [1:0]    _zz_io_result_912;
  wire                _zz_io_result_913;
  reg        [1:0]    _zz_io_result_914;
  wire       [1:0]    _zz_io_result_915;
  reg        [1:0]    _zz_io_result_916;
  wire                _zz_io_result_917;
  reg        [1:0]    _zz_io_result_918;
  wire                _zz_io_result_919;
  reg        [1:0]    _zz_io_result_920;
  wire       [7:0]    _zz_io_result_921;
  reg        [7:0]    _zz_io_result_922;
  reg        [31:0]   _zz_io_result_923;
  wire       [7:0]    _zz_io_result_924;
  reg        [7:0]    _zz_io_result_925;
  wire       [7:0]    _zz_io_result_926;
  reg        [7:0]    _zz_io_result_927;
  wire       [7:0]    _zz_io_result_928;
  reg        [7:0]    _zz_io_result_929;
  wire       [3:0]    _zz_io_result_930;
  wire       [3:0]    _zz_io_result_931;
  wire       [3:0]    _zz_io_result_932;
  reg        [3:0]    _zz_io_result_933;
  reg        [3:0]    _zz_io_result_934;
  wire       [1:0]    _zz_io_result_935;
  wire       [1:0]    _zz_io_result_936;
  wire       [1:0]    _zz_io_result_937;
  wire       [1:0]    _zz_io_result_938;
  wire       [1:0]    _zz_io_result_939;
  wire       [1:0]    _zz_io_result_940;
  wire       [1:0]    _zz_io_result_941;
  wire                _zz_io_result_942;
  reg        [1:0]    _zz_io_result_943;
  wire       [1:0]    _zz_io_result_944;
  reg        [1:0]    _zz_io_result_945;
  wire                _zz_io_result_946;
  reg        [1:0]    _zz_io_result_947;
  wire                _zz_io_result_948;
  reg        [1:0]    _zz_io_result_949;
  wire       [3:0]    _zz_io_result_950;
  wire       [3:0]    _zz_io_result_951;
  reg        [3:0]    _zz_io_result_952;
  wire       [1:0]    _zz_io_result_953;
  wire       [1:0]    _zz_io_result_954;
  wire       [1:0]    _zz_io_result_955;
  reg        [1:0]    _zz_io_result_956;
  wire                _zz_io_result_957;
  reg        [1:0]    _zz_io_result_958;
  wire       [1:0]    _zz_io_result_959;
  wire       [1:0]    _zz_io_result_960;
  reg        [1:0]    _zz_io_result_961;
  wire                _zz_io_result_962;
  reg        [1:0]    _zz_io_result_963;
  wire                _zz_io_result_964;
  reg        [1:0]    _zz_io_result_965;
  reg        [3:0]    _zz_io_result_966;
  wire       [1:0]    _zz_io_result_967;
  wire       [1:0]    _zz_io_result_968;
  wire       [1:0]    _zz_io_result_969;
  wire       [1:0]    _zz_io_result_970;
  wire       [1:0]    _zz_io_result_971;
  wire       [1:0]    _zz_io_result_972;
  wire       [1:0]    _zz_io_result_973;
  wire                _zz_io_result_974;
  reg        [1:0]    _zz_io_result_975;
  wire       [1:0]    _zz_io_result_976;
  reg        [1:0]    _zz_io_result_977;
  wire                _zz_io_result_978;
  reg        [1:0]    _zz_io_result_979;
  wire                _zz_io_result_980;
  reg        [1:0]    _zz_io_result_981;
  reg        [3:0]    _zz_io_result_982;
  wire       [1:0]    _zz_io_result_983;
  wire       [1:0]    _zz_io_result_984;
  wire       [1:0]    _zz_io_result_985;
  wire       [1:0]    _zz_io_result_986;
  wire       [1:0]    _zz_io_result_987;
  wire       [1:0]    _zz_io_result_988;
  wire       [1:0]    _zz_io_result_989;
  wire                _zz_io_result_990;
  reg        [1:0]    _zz_io_result_991;
  wire       [1:0]    _zz_io_result_992;
  reg        [1:0]    _zz_io_result_993;
  wire                _zz_io_result_994;
  reg        [1:0]    _zz_io_result_995;
  wire                _zz_io_result_996;
  reg        [1:0]    _zz_io_result_997;
  wire       [7:0]    _zz_io_result_998;
  reg        [7:0]    _zz_io_result_999;
  wire       [7:0]    _zz_io_result_1000;
  reg        [7:0]    _zz_io_result_1001;
  wire       [7:0]    _zz_io_result_1002;
  reg        [7:0]    _zz_io_result_1003;
  wire       [7:0]    _zz_io_result_1004;
  reg        [7:0]    _zz_io_result_1005;
  wire       [3:0]    _zz_io_result_1006;
  wire       [3:0]    _zz_io_result_1007;
  wire       [3:0]    _zz_io_result_1008;
  reg        [3:0]    _zz_io_result_1009;
  reg        [3:0]    _zz_io_result_1010;
  wire       [1:0]    _zz_io_result_1011;
  wire       [1:0]    _zz_io_result_1012;
  wire       [1:0]    _zz_io_result_1013;
  wire       [1:0]    _zz_io_result_1014;
  wire       [1:0]    _zz_io_result_1015;
  wire       [1:0]    _zz_io_result_1016;
  wire       [1:0]    _zz_io_result_1017;
  wire                _zz_io_result_1018;
  reg        [1:0]    _zz_io_result_1019;
  wire       [1:0]    _zz_io_result_1020;
  reg        [1:0]    _zz_io_result_1021;
  wire                _zz_io_result_1022;
  reg        [1:0]    _zz_io_result_1023;
  wire                _zz_io_result_1024;
  reg        [1:0]    _zz_io_result_1025;
  wire       [3:0]    _zz_io_result_1026;
  wire       [3:0]    _zz_io_result_1027;
  reg        [3:0]    _zz_io_result_1028;
  wire       [1:0]    _zz_io_result_1029;
  wire       [1:0]    _zz_io_result_1030;
  wire       [1:0]    _zz_io_result_1031;
  reg        [1:0]    _zz_io_result_1032;
  wire                _zz_io_result_1033;
  reg        [1:0]    _zz_io_result_1034;
  wire       [1:0]    _zz_io_result_1035;
  wire       [1:0]    _zz_io_result_1036;
  reg        [1:0]    _zz_io_result_1037;
  wire                _zz_io_result_1038;
  reg        [1:0]    _zz_io_result_1039;
  wire                _zz_io_result_1040;
  reg        [1:0]    _zz_io_result_1041;
  reg        [3:0]    _zz_io_result_1042;
  wire       [1:0]    _zz_io_result_1043;
  wire       [1:0]    _zz_io_result_1044;
  wire       [1:0]    _zz_io_result_1045;
  wire       [1:0]    _zz_io_result_1046;
  wire       [1:0]    _zz_io_result_1047;
  wire       [1:0]    _zz_io_result_1048;
  wire       [1:0]    _zz_io_result_1049;
  wire                _zz_io_result_1050;
  reg        [1:0]    _zz_io_result_1051;
  wire       [1:0]    _zz_io_result_1052;
  reg        [1:0]    _zz_io_result_1053;
  wire                _zz_io_result_1054;
  reg        [1:0]    _zz_io_result_1055;
  wire                _zz_io_result_1056;
  reg        [1:0]    _zz_io_result_1057;
  reg        [3:0]    _zz_io_result_1058;
  wire       [1:0]    _zz_io_result_1059;
  wire       [1:0]    _zz_io_result_1060;
  wire       [1:0]    _zz_io_result_1061;
  wire       [1:0]    _zz_io_result_1062;
  wire       [1:0]    _zz_io_result_1063;
  wire       [1:0]    _zz_io_result_1064;
  wire       [1:0]    _zz_io_result_1065;
  wire                _zz_io_result_1066;
  reg        [1:0]    _zz_io_result_1067;
  wire       [1:0]    _zz_io_result_1068;
  reg        [1:0]    _zz_io_result_1069;
  wire                _zz_io_result_1070;
  reg        [1:0]    _zz_io_result_1071;
  wire                _zz_io_result_1072;
  reg        [1:0]    _zz_io_result_1073;
  wire       [7:0]    _zz_io_result_1074;
  reg        [7:0]    _zz_io_result_1075;
  wire       [7:0]    _zz_io_result_1076;
  reg        [7:0]    _zz_io_result_1077;
  wire       [7:0]    _zz_io_result_1078;
  reg        [7:0]    _zz_io_result_1079;
  wire       [7:0]    _zz_io_result_1080;
  reg        [7:0]    _zz_io_result_1081;
  wire       [3:0]    _zz_io_result_1082;
  wire       [3:0]    _zz_io_result_1083;
  wire       [3:0]    _zz_io_result_1084;
  reg        [3:0]    _zz_io_result_1085;
  reg        [3:0]    _zz_io_result_1086;
  wire       [1:0]    _zz_io_result_1087;
  wire       [1:0]    _zz_io_result_1088;
  wire       [1:0]    _zz_io_result_1089;
  wire       [1:0]    _zz_io_result_1090;
  wire       [1:0]    _zz_io_result_1091;
  wire       [1:0]    _zz_io_result_1092;
  wire       [1:0]    _zz_io_result_1093;
  wire                _zz_io_result_1094;
  reg        [1:0]    _zz_io_result_1095;
  wire       [1:0]    _zz_io_result_1096;
  reg        [1:0]    _zz_io_result_1097;
  wire                _zz_io_result_1098;
  reg        [1:0]    _zz_io_result_1099;
  wire                _zz_io_result_1100;
  reg        [1:0]    _zz_io_result_1101;
  wire       [3:0]    _zz_io_result_1102;
  wire       [3:0]    _zz_io_result_1103;
  reg        [3:0]    _zz_io_result_1104;
  wire       [1:0]    _zz_io_result_1105;
  wire       [1:0]    _zz_io_result_1106;
  wire       [1:0]    _zz_io_result_1107;
  reg        [1:0]    _zz_io_result_1108;
  wire                _zz_io_result_1109;
  reg        [1:0]    _zz_io_result_1110;
  wire       [1:0]    _zz_io_result_1111;
  wire       [1:0]    _zz_io_result_1112;
  reg        [1:0]    _zz_io_result_1113;
  wire                _zz_io_result_1114;
  reg        [1:0]    _zz_io_result_1115;
  wire                _zz_io_result_1116;
  reg        [1:0]    _zz_io_result_1117;
  reg        [3:0]    _zz_io_result_1118;
  wire       [1:0]    _zz_io_result_1119;
  wire       [1:0]    _zz_io_result_1120;
  wire       [1:0]    _zz_io_result_1121;
  wire       [1:0]    _zz_io_result_1122;
  wire       [1:0]    _zz_io_result_1123;
  wire       [1:0]    _zz_io_result_1124;
  wire       [1:0]    _zz_io_result_1125;
  wire                _zz_io_result_1126;
  reg        [1:0]    _zz_io_result_1127;
  wire       [1:0]    _zz_io_result_1128;
  reg        [1:0]    _zz_io_result_1129;
  wire                _zz_io_result_1130;
  reg        [1:0]    _zz_io_result_1131;
  wire                _zz_io_result_1132;
  reg        [1:0]    _zz_io_result_1133;
  reg        [3:0]    _zz_io_result_1134;
  wire       [1:0]    _zz_io_result_1135;
  wire       [1:0]    _zz_io_result_1136;
  wire       [1:0]    _zz_io_result_1137;
  wire       [1:0]    _zz_io_result_1138;
  wire       [1:0]    _zz_io_result_1139;
  wire       [1:0]    _zz_io_result_1140;
  wire       [1:0]    _zz_io_result_1141;
  wire                _zz_io_result_1142;
  reg        [1:0]    _zz_io_result_1143;
  wire       [1:0]    _zz_io_result_1144;
  reg        [1:0]    _zz_io_result_1145;
  wire                _zz_io_result_1146;
  reg        [1:0]    _zz_io_result_1147;
  wire                _zz_io_result_1148;
  reg        [1:0]    _zz_io_result_1149;
  wire       [7:0]    _zz_io_result_1150;
  reg        [7:0]    _zz_io_result_1151;
  wire       [7:0]    _zz_io_result_1152;
  reg        [7:0]    _zz_io_result_1153;
  wire       [7:0]    _zz_io_result_1154;
  reg        [7:0]    _zz_io_result_1155;
  wire       [7:0]    _zz_io_result_1156;
  reg        [7:0]    _zz_io_result_1157;
  wire       [3:0]    _zz_io_result_1158;
  wire       [3:0]    _zz_io_result_1159;
  wire       [3:0]    _zz_io_result_1160;
  reg        [3:0]    _zz_io_result_1161;
  reg        [3:0]    _zz_io_result_1162;
  wire       [1:0]    _zz_io_result_1163;
  wire       [1:0]    _zz_io_result_1164;
  wire       [1:0]    _zz_io_result_1165;
  wire       [1:0]    _zz_io_result_1166;
  wire       [1:0]    _zz_io_result_1167;
  wire       [1:0]    _zz_io_result_1168;
  wire       [1:0]    _zz_io_result_1169;
  wire                _zz_io_result_1170;
  reg        [1:0]    _zz_io_result_1171;
  wire       [1:0]    _zz_io_result_1172;
  reg        [1:0]    _zz_io_result_1173;
  wire                _zz_io_result_1174;
  reg        [1:0]    _zz_io_result_1175;
  wire                _zz_io_result_1176;
  reg        [1:0]    _zz_io_result_1177;
  wire       [3:0]    _zz_io_result_1178;
  wire       [3:0]    _zz_io_result_1179;
  reg        [3:0]    _zz_io_result_1180;
  wire       [1:0]    _zz_io_result_1181;
  wire       [1:0]    _zz_io_result_1182;
  wire       [1:0]    _zz_io_result_1183;
  reg        [1:0]    _zz_io_result_1184;
  wire                _zz_io_result_1185;
  reg        [1:0]    _zz_io_result_1186;
  wire       [1:0]    _zz_io_result_1187;
  wire       [1:0]    _zz_io_result_1188;
  reg        [1:0]    _zz_io_result_1189;
  wire                _zz_io_result_1190;
  reg        [1:0]    _zz_io_result_1191;
  wire                _zz_io_result_1192;
  reg        [1:0]    _zz_io_result_1193;
  reg        [3:0]    _zz_io_result_1194;
  wire       [1:0]    _zz_io_result_1195;
  wire       [1:0]    _zz_io_result_1196;
  wire       [1:0]    _zz_io_result_1197;
  wire       [1:0]    _zz_io_result_1198;
  wire       [1:0]    _zz_io_result_1199;
  wire       [1:0]    _zz_io_result_1200;
  wire       [1:0]    _zz_io_result_1201;
  wire                _zz_io_result_1202;
  reg        [1:0]    _zz_io_result_1203;
  wire       [1:0]    _zz_io_result_1204;
  reg        [1:0]    _zz_io_result_1205;
  wire                _zz_io_result_1206;
  reg        [1:0]    _zz_io_result_1207;
  wire                _zz_io_result_1208;
  reg        [1:0]    _zz_io_result_1209;
  reg        [3:0]    _zz_io_result_1210;
  wire       [1:0]    _zz_io_result_1211;
  wire       [1:0]    _zz_io_result_1212;
  wire       [1:0]    _zz_io_result_1213;
  wire       [1:0]    _zz_io_result_1214;
  wire       [1:0]    _zz_io_result_1215;
  wire       [1:0]    _zz_io_result_1216;
  wire       [1:0]    _zz_io_result_1217;
  wire                _zz_io_result_1218;
  reg        [1:0]    _zz_io_result_1219;
  wire       [1:0]    _zz_io_result_1220;
  reg        [1:0]    _zz_io_result_1221;
  wire                _zz_io_result_1222;
  reg        [1:0]    _zz_io_result_1223;
  wire                _zz_io_result_1224;
  reg        [1:0]    _zz_io_result_1225;
  wire       [7:0]    _zz_io_result_1226;
  reg        [7:0]    _zz_io_result_1227;
  wire       [127:0]  _zz_io_result_1228;
  wire       [31:0]   _zz_io_result_1229;
  wire       [31:0]   _zz_io_result_1230;
  wire       [31:0]   _zz_io_result_1231;
  wire       [31:0]   _zz_io_result_1232;
  wire       [127:0]  _zz_io_result_1233;
  reg        [31:0]   _zz_io_result_1234;
  wire       [31:0]   _zz_io_result_1235;
  wire       [7:0]    _zz_io_result_1236;
  wire       [7:0]    _zz_io_result_1237;
  reg        [7:0]    _zz_io_result_1238;
  wire       [31:0]   _zz_io_result_1239;
  wire       [7:0]    _zz_io_result_1240;
  wire       [7:0]    _zz_io_result_1241;
  reg        [7:0]    _zz_io_result_1242;
  wire       [31:0]   _zz_io_result_1243;
  wire       [7:0]    _zz_io_result_1244;
  wire       [7:0]    _zz_io_result_1245;
  reg        [7:0]    _zz_io_result_1246;
  wire       [31:0]   _zz_io_result_1247;
  wire       [7:0]    _zz_io_result_1248;
  wire       [7:0]    _zz_io_result_1249;
  reg        [7:0]    _zz_io_result_1250;
  reg        [31:0]   _zz_io_result_1251;
  wire       [31:0]   _zz_io_result_1252;
  wire       [7:0]    _zz_io_result_1253;
  wire       [7:0]    _zz_io_result_1254;
  reg        [7:0]    _zz_io_result_1255;
  wire       [31:0]   _zz_io_result_1256;
  wire       [7:0]    _zz_io_result_1257;
  wire       [7:0]    _zz_io_result_1258;
  reg        [7:0]    _zz_io_result_1259;
  wire       [31:0]   _zz_io_result_1260;
  wire       [7:0]    _zz_io_result_1261;
  wire       [7:0]    _zz_io_result_1262;
  reg        [7:0]    _zz_io_result_1263;
  wire       [31:0]   _zz_io_result_1264;
  wire       [7:0]    _zz_io_result_1265;
  wire       [7:0]    _zz_io_result_1266;
  reg        [7:0]    _zz_io_result_1267;
  reg        [31:0]   _zz_io_result_1268;
  wire       [31:0]   _zz_io_result_1269;
  wire       [7:0]    _zz_io_result_1270;
  wire       [7:0]    _zz_io_result_1271;
  reg        [7:0]    _zz_io_result_1272;
  wire       [31:0]   _zz_io_result_1273;
  wire       [7:0]    _zz_io_result_1274;
  wire       [7:0]    _zz_io_result_1275;
  reg        [7:0]    _zz_io_result_1276;
  wire       [31:0]   _zz_io_result_1277;
  wire       [7:0]    _zz_io_result_1278;
  wire       [7:0]    _zz_io_result_1279;
  reg        [7:0]    _zz_io_result_1280;
  wire       [31:0]   _zz_io_result_1281;
  wire       [7:0]    _zz_io_result_1282;
  wire       [7:0]    _zz_io_result_1283;
  reg        [7:0]    _zz_io_result_1284;
  reg        [31:0]   _zz_io_result_1285;
  wire       [31:0]   _zz_io_result_1286;
  wire       [7:0]    _zz_io_result_1287;
  wire       [7:0]    _zz_io_result_1288;
  reg        [7:0]    _zz_io_result_1289;
  wire       [31:0]   _zz_io_result_1290;
  wire       [7:0]    _zz_io_result_1291;
  wire       [7:0]    _zz_io_result_1292;
  reg        [7:0]    _zz_io_result_1293;
  wire       [31:0]   _zz_io_result_1294;
  wire       [7:0]    _zz_io_result_1295;
  wire       [7:0]    _zz_io_result_1296;
  reg        [7:0]    _zz_io_result_1297;
  wire       [31:0]   _zz_io_result_1298;
  wire       [7:0]    _zz_io_result_1299;
  wire       [7:0]    _zz_io_result_1300;
  reg        [7:0]    _zz_io_result_1301;

  assign _zz_io_result = io_roundData[31 : 0];
  assign _zz_io_result_1 = io_roundData[63 : 32];
  assign _zz_io_result_2 = io_roundData[95 : 64];
  assign _zz_io_result_3 = io_roundData[127 : 96];
  assign _zz_io_result_9 = _zz_io_result[7 : 0];
  always @(*) begin
    _zz_io_result_12[7] = (((((_zz_io_result_9[7] ^ _zz_io_result_9[6]) ^ _zz_io_result_9[5]) ^ _zz_io_result_9[2]) ^ _zz_io_result_9[1]) ^ _zz_io_result_9[0]);
    _zz_io_result_12[6] = (((_zz_io_result_9[6] ^ _zz_io_result_9[5]) ^ _zz_io_result_9[4]) ^ _zz_io_result_9[0]);
    _zz_io_result_12[5] = (((_zz_io_result_9[6] ^ _zz_io_result_9[5]) ^ _zz_io_result_9[1]) ^ _zz_io_result_9[0]);
    _zz_io_result_12[4] = (((_zz_io_result_9[7] ^ _zz_io_result_9[6]) ^ _zz_io_result_9[5]) ^ _zz_io_result_9[0]);
    _zz_io_result_12[3] = ((((_zz_io_result_9[7] ^ _zz_io_result_9[4]) ^ _zz_io_result_9[3]) ^ _zz_io_result_9[1]) ^ _zz_io_result_9[0]);
    _zz_io_result_12[2] = _zz_io_result_9[0];
    _zz_io_result_12[1] = ((_zz_io_result_9[6] ^ _zz_io_result_9[5]) ^ _zz_io_result_9[0]);
    _zz_io_result_12[0] = ((((_zz_io_result_9[6] ^ _zz_io_result_9[3]) ^ _zz_io_result_9[2]) ^ _zz_io_result_9[1]) ^ _zz_io_result_9[0]);
  end

  assign _zz_io_result_11 = _zz_io_result_12;
  assign _zz_io_result_15 = _zz_io_result_11[7 : 4];
  assign _zz_io_result_16 = _zz_io_result_11[3 : 0];
  assign _zz_io_result_17 = (_zz_io_result_15 ^ _zz_io_result_16);
  always @(*) begin
    _zz_io_result_18[3] = (_zz_io_result_17[2] ^ _zz_io_result_17[0]);
    _zz_io_result_18[2] = (_zz_io_result_17[3] ^ _zz_io_result_17[1]);
    _zz_io_result_18[1] = (_zz_io_result_17[1] ^ _zz_io_result_17[0]);
    _zz_io_result_18[0] = _zz_io_result_17[0];
  end

  assign _zz_io_result_20 = _zz_io_result_15[3 : 2];
  assign _zz_io_result_21 = _zz_io_result_15[1 : 0];
  assign _zz_io_result_22 = _zz_io_result_16[3 : 2];
  assign _zz_io_result_23 = _zz_io_result_16[1 : 0];
  assign _zz_io_result_24 = (_zz_io_result_20 ^ _zz_io_result_21);
  assign _zz_io_result_25 = (_zz_io_result_22 ^ _zz_io_result_23);
  assign _zz_io_result_27 = ((_zz_io_result_25[0] && _zz_io_result_24[1]) ^ (_zz_io_result_24[0] && _zz_io_result_25[1]));
  always @(*) begin
    _zz_io_result_28[1] = ((_zz_io_result_25[0] && _zz_io_result_24[0]) ^ _zz_io_result_27);
    _zz_io_result_28[0] = ((_zz_io_result_25[1] && _zz_io_result_24[1]) ^ _zz_io_result_27);
  end

  assign _zz_io_result_26 = _zz_io_result_28;
  always @(*) begin
    _zz_io_result_30[1] = _zz_io_result_26[0];
    _zz_io_result_30[0] = (_zz_io_result_26[0] ^ _zz_io_result_26[1]);
  end

  assign _zz_io_result_29 = _zz_io_result_30;
  assign _zz_io_result_31 = ((_zz_io_result_22[0] && _zz_io_result_20[1]) ^ (_zz_io_result_20[0] && _zz_io_result_22[1]));
  always @(*) begin
    _zz_io_result_32[1] = ((_zz_io_result_22[0] && _zz_io_result_20[0]) ^ _zz_io_result_31);
    _zz_io_result_32[0] = ((_zz_io_result_22[1] && _zz_io_result_20[1]) ^ _zz_io_result_31);
  end

  assign _zz_io_result_33 = ((_zz_io_result_23[0] && _zz_io_result_21[1]) ^ (_zz_io_result_21[0] && _zz_io_result_23[1]));
  always @(*) begin
    _zz_io_result_34[1] = ((_zz_io_result_23[0] && _zz_io_result_21[0]) ^ _zz_io_result_33);
    _zz_io_result_34[0] = ((_zz_io_result_23[1] && _zz_io_result_21[1]) ^ _zz_io_result_33);
  end

  always @(*) begin
    _zz_io_result_19[3 : 2] = (_zz_io_result_32 ^ _zz_io_result_29);
    _zz_io_result_19[1 : 0] = (_zz_io_result_34 ^ _zz_io_result_29);
  end

  assign _zz_io_result_35 = (_zz_io_result_18 ^ _zz_io_result_19);
  assign _zz_io_result_38 = _zz_io_result_35[3 : 2];
  assign _zz_io_result_39 = _zz_io_result_35[1 : 0];
  assign _zz_io_result_40 = (_zz_io_result_38 ^ _zz_io_result_39);
  always @(*) begin
    _zz_io_result_41[1] = _zz_io_result_40[1];
    _zz_io_result_41[0] = (_zz_io_result_40[0] ^ _zz_io_result_40[1]);
  end

  assign _zz_io_result_42 = ((_zz_io_result_39[0] && _zz_io_result_38[1]) ^ (_zz_io_result_38[0] && _zz_io_result_39[1]));
  always @(*) begin
    _zz_io_result_43[1] = ((_zz_io_result_39[0] && _zz_io_result_38[0]) ^ _zz_io_result_42);
    _zz_io_result_43[0] = ((_zz_io_result_39[1] && _zz_io_result_38[1]) ^ _zz_io_result_42);
  end

  assign _zz_io_result_44 = (_zz_io_result_41 ^ _zz_io_result_43);
  always @(*) begin
    _zz_io_result_46[1] = _zz_io_result_44[0];
    _zz_io_result_46[0] = _zz_io_result_44[1];
  end

  assign _zz_io_result_45 = _zz_io_result_46;
  assign _zz_io_result_47 = ((_zz_io_result_45[0] && _zz_io_result_38[1]) ^ (_zz_io_result_38[0] && _zz_io_result_45[1]));
  always @(*) begin
    _zz_io_result_48[1] = ((_zz_io_result_45[0] && _zz_io_result_38[0]) ^ _zz_io_result_47);
    _zz_io_result_48[0] = ((_zz_io_result_45[1] && _zz_io_result_38[1]) ^ _zz_io_result_47);
  end

  assign _zz_io_result_49 = ((_zz_io_result_45[0] && _zz_io_result_39[1]) ^ (_zz_io_result_39[0] && _zz_io_result_45[1]));
  always @(*) begin
    _zz_io_result_50[1] = ((_zz_io_result_45[0] && _zz_io_result_39[0]) ^ _zz_io_result_49);
    _zz_io_result_50[0] = ((_zz_io_result_45[1] && _zz_io_result_39[1]) ^ _zz_io_result_49);
  end

  always @(*) begin
    _zz_io_result_37[3 : 2] = _zz_io_result_50;
    _zz_io_result_37[1 : 0] = _zz_io_result_48;
  end

  assign _zz_io_result_36 = _zz_io_result_37;
  assign _zz_io_result_52 = _zz_io_result_15[3 : 2];
  assign _zz_io_result_53 = _zz_io_result_15[1 : 0];
  assign _zz_io_result_54 = _zz_io_result_36[3 : 2];
  assign _zz_io_result_55 = _zz_io_result_36[1 : 0];
  assign _zz_io_result_56 = (_zz_io_result_52 ^ _zz_io_result_53);
  assign _zz_io_result_57 = (_zz_io_result_54 ^ _zz_io_result_55);
  assign _zz_io_result_59 = ((_zz_io_result_57[0] && _zz_io_result_56[1]) ^ (_zz_io_result_56[0] && _zz_io_result_57[1]));
  always @(*) begin
    _zz_io_result_60[1] = ((_zz_io_result_57[0] && _zz_io_result_56[0]) ^ _zz_io_result_59);
    _zz_io_result_60[0] = ((_zz_io_result_57[1] && _zz_io_result_56[1]) ^ _zz_io_result_59);
  end

  assign _zz_io_result_58 = _zz_io_result_60;
  always @(*) begin
    _zz_io_result_62[1] = _zz_io_result_58[0];
    _zz_io_result_62[0] = (_zz_io_result_58[0] ^ _zz_io_result_58[1]);
  end

  assign _zz_io_result_61 = _zz_io_result_62;
  assign _zz_io_result_63 = ((_zz_io_result_54[0] && _zz_io_result_52[1]) ^ (_zz_io_result_52[0] && _zz_io_result_54[1]));
  always @(*) begin
    _zz_io_result_64[1] = ((_zz_io_result_54[0] && _zz_io_result_52[0]) ^ _zz_io_result_63);
    _zz_io_result_64[0] = ((_zz_io_result_54[1] && _zz_io_result_52[1]) ^ _zz_io_result_63);
  end

  assign _zz_io_result_65 = ((_zz_io_result_55[0] && _zz_io_result_53[1]) ^ (_zz_io_result_53[0] && _zz_io_result_55[1]));
  always @(*) begin
    _zz_io_result_66[1] = ((_zz_io_result_55[0] && _zz_io_result_53[0]) ^ _zz_io_result_65);
    _zz_io_result_66[0] = ((_zz_io_result_55[1] && _zz_io_result_53[1]) ^ _zz_io_result_65);
  end

  always @(*) begin
    _zz_io_result_51[3 : 2] = (_zz_io_result_64 ^ _zz_io_result_61);
    _zz_io_result_51[1 : 0] = (_zz_io_result_66 ^ _zz_io_result_61);
  end

  assign _zz_io_result_68 = _zz_io_result_16[3 : 2];
  assign _zz_io_result_69 = _zz_io_result_16[1 : 0];
  assign _zz_io_result_70 = _zz_io_result_36[3 : 2];
  assign _zz_io_result_71 = _zz_io_result_36[1 : 0];
  assign _zz_io_result_72 = (_zz_io_result_68 ^ _zz_io_result_69);
  assign _zz_io_result_73 = (_zz_io_result_70 ^ _zz_io_result_71);
  assign _zz_io_result_75 = ((_zz_io_result_73[0] && _zz_io_result_72[1]) ^ (_zz_io_result_72[0] && _zz_io_result_73[1]));
  always @(*) begin
    _zz_io_result_76[1] = ((_zz_io_result_73[0] && _zz_io_result_72[0]) ^ _zz_io_result_75);
    _zz_io_result_76[0] = ((_zz_io_result_73[1] && _zz_io_result_72[1]) ^ _zz_io_result_75);
  end

  assign _zz_io_result_74 = _zz_io_result_76;
  always @(*) begin
    _zz_io_result_78[1] = _zz_io_result_74[0];
    _zz_io_result_78[0] = (_zz_io_result_74[0] ^ _zz_io_result_74[1]);
  end

  assign _zz_io_result_77 = _zz_io_result_78;
  assign _zz_io_result_79 = ((_zz_io_result_70[0] && _zz_io_result_68[1]) ^ (_zz_io_result_68[0] && _zz_io_result_70[1]));
  always @(*) begin
    _zz_io_result_80[1] = ((_zz_io_result_70[0] && _zz_io_result_68[0]) ^ _zz_io_result_79);
    _zz_io_result_80[0] = ((_zz_io_result_70[1] && _zz_io_result_68[1]) ^ _zz_io_result_79);
  end

  assign _zz_io_result_81 = ((_zz_io_result_71[0] && _zz_io_result_69[1]) ^ (_zz_io_result_69[0] && _zz_io_result_71[1]));
  always @(*) begin
    _zz_io_result_82[1] = ((_zz_io_result_71[0] && _zz_io_result_69[0]) ^ _zz_io_result_81);
    _zz_io_result_82[0] = ((_zz_io_result_71[1] && _zz_io_result_69[1]) ^ _zz_io_result_81);
  end

  always @(*) begin
    _zz_io_result_67[3 : 2] = (_zz_io_result_80 ^ _zz_io_result_77);
    _zz_io_result_67[1 : 0] = (_zz_io_result_82 ^ _zz_io_result_77);
  end

  always @(*) begin
    _zz_io_result_14[7 : 4] = _zz_io_result_67;
    _zz_io_result_14[3 : 0] = _zz_io_result_51;
  end

  assign _zz_io_result_13 = _zz_io_result_14;
  always @(*) begin
    _zz_io_result_84[7] = (_zz_io_result_13[5] ^ _zz_io_result_13[3]);
    _zz_io_result_84[6] = (_zz_io_result_13[7] ^ _zz_io_result_13[3]);
    _zz_io_result_84[5] = (_zz_io_result_13[6] ^ _zz_io_result_13[0]);
    _zz_io_result_84[4] = ((_zz_io_result_13[7] ^ _zz_io_result_13[5]) ^ _zz_io_result_13[3]);
    _zz_io_result_84[3] = ((((_zz_io_result_13[7] ^ _zz_io_result_13[6]) ^ _zz_io_result_13[5]) ^ _zz_io_result_13[4]) ^ _zz_io_result_13[3]);
    _zz_io_result_84[2] = ((((_zz_io_result_13[6] ^ _zz_io_result_13[5]) ^ _zz_io_result_13[3]) ^ _zz_io_result_13[2]) ^ _zz_io_result_13[0]);
    _zz_io_result_84[1] = ((_zz_io_result_13[5] ^ _zz_io_result_13[4]) ^ _zz_io_result_13[1]);
    _zz_io_result_84[0] = ((_zz_io_result_13[6] ^ _zz_io_result_13[4]) ^ _zz_io_result_13[1]);
  end

  assign _zz_io_result_83 = _zz_io_result_84;
  always @(*) begin
    _zz_io_result_10[7] = _zz_io_result_83[7];
    _zz_io_result_10[6] = (! _zz_io_result_83[6]);
    _zz_io_result_10[5] = (! _zz_io_result_83[5]);
    _zz_io_result_10[4] = _zz_io_result_83[4];
    _zz_io_result_10[3] = _zz_io_result_83[3];
    _zz_io_result_10[2] = _zz_io_result_83[2];
    _zz_io_result_10[1] = (! _zz_io_result_83[1]);
    _zz_io_result_10[0] = (! _zz_io_result_83[0]);
  end

  always @(*) begin
    _zz_io_result_8[7 : 0] = _zz_io_result_10;
    _zz_io_result_8[15 : 8] = _zz_io_result_86;
    _zz_io_result_8[23 : 16] = _zz_io_result_162;
    _zz_io_result_8[31 : 24] = _zz_io_result_238;
  end

  assign _zz_io_result_85 = _zz_io_result[15 : 8];
  always @(*) begin
    _zz_io_result_88[7] = (((((_zz_io_result_85[7] ^ _zz_io_result_85[6]) ^ _zz_io_result_85[5]) ^ _zz_io_result_85[2]) ^ _zz_io_result_85[1]) ^ _zz_io_result_85[0]);
    _zz_io_result_88[6] = (((_zz_io_result_85[6] ^ _zz_io_result_85[5]) ^ _zz_io_result_85[4]) ^ _zz_io_result_85[0]);
    _zz_io_result_88[5] = (((_zz_io_result_85[6] ^ _zz_io_result_85[5]) ^ _zz_io_result_85[1]) ^ _zz_io_result_85[0]);
    _zz_io_result_88[4] = (((_zz_io_result_85[7] ^ _zz_io_result_85[6]) ^ _zz_io_result_85[5]) ^ _zz_io_result_85[0]);
    _zz_io_result_88[3] = ((((_zz_io_result_85[7] ^ _zz_io_result_85[4]) ^ _zz_io_result_85[3]) ^ _zz_io_result_85[1]) ^ _zz_io_result_85[0]);
    _zz_io_result_88[2] = _zz_io_result_85[0];
    _zz_io_result_88[1] = ((_zz_io_result_85[6] ^ _zz_io_result_85[5]) ^ _zz_io_result_85[0]);
    _zz_io_result_88[0] = ((((_zz_io_result_85[6] ^ _zz_io_result_85[3]) ^ _zz_io_result_85[2]) ^ _zz_io_result_85[1]) ^ _zz_io_result_85[0]);
  end

  assign _zz_io_result_87 = _zz_io_result_88;
  assign _zz_io_result_91 = _zz_io_result_87[7 : 4];
  assign _zz_io_result_92 = _zz_io_result_87[3 : 0];
  assign _zz_io_result_93 = (_zz_io_result_91 ^ _zz_io_result_92);
  always @(*) begin
    _zz_io_result_94[3] = (_zz_io_result_93[2] ^ _zz_io_result_93[0]);
    _zz_io_result_94[2] = (_zz_io_result_93[3] ^ _zz_io_result_93[1]);
    _zz_io_result_94[1] = (_zz_io_result_93[1] ^ _zz_io_result_93[0]);
    _zz_io_result_94[0] = _zz_io_result_93[0];
  end

  assign _zz_io_result_96 = _zz_io_result_91[3 : 2];
  assign _zz_io_result_97 = _zz_io_result_91[1 : 0];
  assign _zz_io_result_98 = _zz_io_result_92[3 : 2];
  assign _zz_io_result_99 = _zz_io_result_92[1 : 0];
  assign _zz_io_result_100 = (_zz_io_result_96 ^ _zz_io_result_97);
  assign _zz_io_result_101 = (_zz_io_result_98 ^ _zz_io_result_99);
  assign _zz_io_result_103 = ((_zz_io_result_101[0] && _zz_io_result_100[1]) ^ (_zz_io_result_100[0] && _zz_io_result_101[1]));
  always @(*) begin
    _zz_io_result_104[1] = ((_zz_io_result_101[0] && _zz_io_result_100[0]) ^ _zz_io_result_103);
    _zz_io_result_104[0] = ((_zz_io_result_101[1] && _zz_io_result_100[1]) ^ _zz_io_result_103);
  end

  assign _zz_io_result_102 = _zz_io_result_104;
  always @(*) begin
    _zz_io_result_106[1] = _zz_io_result_102[0];
    _zz_io_result_106[0] = (_zz_io_result_102[0] ^ _zz_io_result_102[1]);
  end

  assign _zz_io_result_105 = _zz_io_result_106;
  assign _zz_io_result_107 = ((_zz_io_result_98[0] && _zz_io_result_96[1]) ^ (_zz_io_result_96[0] && _zz_io_result_98[1]));
  always @(*) begin
    _zz_io_result_108[1] = ((_zz_io_result_98[0] && _zz_io_result_96[0]) ^ _zz_io_result_107);
    _zz_io_result_108[0] = ((_zz_io_result_98[1] && _zz_io_result_96[1]) ^ _zz_io_result_107);
  end

  assign _zz_io_result_109 = ((_zz_io_result_99[0] && _zz_io_result_97[1]) ^ (_zz_io_result_97[0] && _zz_io_result_99[1]));
  always @(*) begin
    _zz_io_result_110[1] = ((_zz_io_result_99[0] && _zz_io_result_97[0]) ^ _zz_io_result_109);
    _zz_io_result_110[0] = ((_zz_io_result_99[1] && _zz_io_result_97[1]) ^ _zz_io_result_109);
  end

  always @(*) begin
    _zz_io_result_95[3 : 2] = (_zz_io_result_108 ^ _zz_io_result_105);
    _zz_io_result_95[1 : 0] = (_zz_io_result_110 ^ _zz_io_result_105);
  end

  assign _zz_io_result_111 = (_zz_io_result_94 ^ _zz_io_result_95);
  assign _zz_io_result_114 = _zz_io_result_111[3 : 2];
  assign _zz_io_result_115 = _zz_io_result_111[1 : 0];
  assign _zz_io_result_116 = (_zz_io_result_114 ^ _zz_io_result_115);
  always @(*) begin
    _zz_io_result_117[1] = _zz_io_result_116[1];
    _zz_io_result_117[0] = (_zz_io_result_116[0] ^ _zz_io_result_116[1]);
  end

  assign _zz_io_result_118 = ((_zz_io_result_115[0] && _zz_io_result_114[1]) ^ (_zz_io_result_114[0] && _zz_io_result_115[1]));
  always @(*) begin
    _zz_io_result_119[1] = ((_zz_io_result_115[0] && _zz_io_result_114[0]) ^ _zz_io_result_118);
    _zz_io_result_119[0] = ((_zz_io_result_115[1] && _zz_io_result_114[1]) ^ _zz_io_result_118);
  end

  assign _zz_io_result_120 = (_zz_io_result_117 ^ _zz_io_result_119);
  always @(*) begin
    _zz_io_result_122[1] = _zz_io_result_120[0];
    _zz_io_result_122[0] = _zz_io_result_120[1];
  end

  assign _zz_io_result_121 = _zz_io_result_122;
  assign _zz_io_result_123 = ((_zz_io_result_121[0] && _zz_io_result_114[1]) ^ (_zz_io_result_114[0] && _zz_io_result_121[1]));
  always @(*) begin
    _zz_io_result_124[1] = ((_zz_io_result_121[0] && _zz_io_result_114[0]) ^ _zz_io_result_123);
    _zz_io_result_124[0] = ((_zz_io_result_121[1] && _zz_io_result_114[1]) ^ _zz_io_result_123);
  end

  assign _zz_io_result_125 = ((_zz_io_result_121[0] && _zz_io_result_115[1]) ^ (_zz_io_result_115[0] && _zz_io_result_121[1]));
  always @(*) begin
    _zz_io_result_126[1] = ((_zz_io_result_121[0] && _zz_io_result_115[0]) ^ _zz_io_result_125);
    _zz_io_result_126[0] = ((_zz_io_result_121[1] && _zz_io_result_115[1]) ^ _zz_io_result_125);
  end

  always @(*) begin
    _zz_io_result_113[3 : 2] = _zz_io_result_126;
    _zz_io_result_113[1 : 0] = _zz_io_result_124;
  end

  assign _zz_io_result_112 = _zz_io_result_113;
  assign _zz_io_result_128 = _zz_io_result_91[3 : 2];
  assign _zz_io_result_129 = _zz_io_result_91[1 : 0];
  assign _zz_io_result_130 = _zz_io_result_112[3 : 2];
  assign _zz_io_result_131 = _zz_io_result_112[1 : 0];
  assign _zz_io_result_132 = (_zz_io_result_128 ^ _zz_io_result_129);
  assign _zz_io_result_133 = (_zz_io_result_130 ^ _zz_io_result_131);
  assign _zz_io_result_135 = ((_zz_io_result_133[0] && _zz_io_result_132[1]) ^ (_zz_io_result_132[0] && _zz_io_result_133[1]));
  always @(*) begin
    _zz_io_result_136[1] = ((_zz_io_result_133[0] && _zz_io_result_132[0]) ^ _zz_io_result_135);
    _zz_io_result_136[0] = ((_zz_io_result_133[1] && _zz_io_result_132[1]) ^ _zz_io_result_135);
  end

  assign _zz_io_result_134 = _zz_io_result_136;
  always @(*) begin
    _zz_io_result_138[1] = _zz_io_result_134[0];
    _zz_io_result_138[0] = (_zz_io_result_134[0] ^ _zz_io_result_134[1]);
  end

  assign _zz_io_result_137 = _zz_io_result_138;
  assign _zz_io_result_139 = ((_zz_io_result_130[0] && _zz_io_result_128[1]) ^ (_zz_io_result_128[0] && _zz_io_result_130[1]));
  always @(*) begin
    _zz_io_result_140[1] = ((_zz_io_result_130[0] && _zz_io_result_128[0]) ^ _zz_io_result_139);
    _zz_io_result_140[0] = ((_zz_io_result_130[1] && _zz_io_result_128[1]) ^ _zz_io_result_139);
  end

  assign _zz_io_result_141 = ((_zz_io_result_131[0] && _zz_io_result_129[1]) ^ (_zz_io_result_129[0] && _zz_io_result_131[1]));
  always @(*) begin
    _zz_io_result_142[1] = ((_zz_io_result_131[0] && _zz_io_result_129[0]) ^ _zz_io_result_141);
    _zz_io_result_142[0] = ((_zz_io_result_131[1] && _zz_io_result_129[1]) ^ _zz_io_result_141);
  end

  always @(*) begin
    _zz_io_result_127[3 : 2] = (_zz_io_result_140 ^ _zz_io_result_137);
    _zz_io_result_127[1 : 0] = (_zz_io_result_142 ^ _zz_io_result_137);
  end

  assign _zz_io_result_144 = _zz_io_result_92[3 : 2];
  assign _zz_io_result_145 = _zz_io_result_92[1 : 0];
  assign _zz_io_result_146 = _zz_io_result_112[3 : 2];
  assign _zz_io_result_147 = _zz_io_result_112[1 : 0];
  assign _zz_io_result_148 = (_zz_io_result_144 ^ _zz_io_result_145);
  assign _zz_io_result_149 = (_zz_io_result_146 ^ _zz_io_result_147);
  assign _zz_io_result_151 = ((_zz_io_result_149[0] && _zz_io_result_148[1]) ^ (_zz_io_result_148[0] && _zz_io_result_149[1]));
  always @(*) begin
    _zz_io_result_152[1] = ((_zz_io_result_149[0] && _zz_io_result_148[0]) ^ _zz_io_result_151);
    _zz_io_result_152[0] = ((_zz_io_result_149[1] && _zz_io_result_148[1]) ^ _zz_io_result_151);
  end

  assign _zz_io_result_150 = _zz_io_result_152;
  always @(*) begin
    _zz_io_result_154[1] = _zz_io_result_150[0];
    _zz_io_result_154[0] = (_zz_io_result_150[0] ^ _zz_io_result_150[1]);
  end

  assign _zz_io_result_153 = _zz_io_result_154;
  assign _zz_io_result_155 = ((_zz_io_result_146[0] && _zz_io_result_144[1]) ^ (_zz_io_result_144[0] && _zz_io_result_146[1]));
  always @(*) begin
    _zz_io_result_156[1] = ((_zz_io_result_146[0] && _zz_io_result_144[0]) ^ _zz_io_result_155);
    _zz_io_result_156[0] = ((_zz_io_result_146[1] && _zz_io_result_144[1]) ^ _zz_io_result_155);
  end

  assign _zz_io_result_157 = ((_zz_io_result_147[0] && _zz_io_result_145[1]) ^ (_zz_io_result_145[0] && _zz_io_result_147[1]));
  always @(*) begin
    _zz_io_result_158[1] = ((_zz_io_result_147[0] && _zz_io_result_145[0]) ^ _zz_io_result_157);
    _zz_io_result_158[0] = ((_zz_io_result_147[1] && _zz_io_result_145[1]) ^ _zz_io_result_157);
  end

  always @(*) begin
    _zz_io_result_143[3 : 2] = (_zz_io_result_156 ^ _zz_io_result_153);
    _zz_io_result_143[1 : 0] = (_zz_io_result_158 ^ _zz_io_result_153);
  end

  always @(*) begin
    _zz_io_result_90[7 : 4] = _zz_io_result_143;
    _zz_io_result_90[3 : 0] = _zz_io_result_127;
  end

  assign _zz_io_result_89 = _zz_io_result_90;
  always @(*) begin
    _zz_io_result_160[7] = (_zz_io_result_89[5] ^ _zz_io_result_89[3]);
    _zz_io_result_160[6] = (_zz_io_result_89[7] ^ _zz_io_result_89[3]);
    _zz_io_result_160[5] = (_zz_io_result_89[6] ^ _zz_io_result_89[0]);
    _zz_io_result_160[4] = ((_zz_io_result_89[7] ^ _zz_io_result_89[5]) ^ _zz_io_result_89[3]);
    _zz_io_result_160[3] = ((((_zz_io_result_89[7] ^ _zz_io_result_89[6]) ^ _zz_io_result_89[5]) ^ _zz_io_result_89[4]) ^ _zz_io_result_89[3]);
    _zz_io_result_160[2] = ((((_zz_io_result_89[6] ^ _zz_io_result_89[5]) ^ _zz_io_result_89[3]) ^ _zz_io_result_89[2]) ^ _zz_io_result_89[0]);
    _zz_io_result_160[1] = ((_zz_io_result_89[5] ^ _zz_io_result_89[4]) ^ _zz_io_result_89[1]);
    _zz_io_result_160[0] = ((_zz_io_result_89[6] ^ _zz_io_result_89[4]) ^ _zz_io_result_89[1]);
  end

  assign _zz_io_result_159 = _zz_io_result_160;
  always @(*) begin
    _zz_io_result_86[7] = _zz_io_result_159[7];
    _zz_io_result_86[6] = (! _zz_io_result_159[6]);
    _zz_io_result_86[5] = (! _zz_io_result_159[5]);
    _zz_io_result_86[4] = _zz_io_result_159[4];
    _zz_io_result_86[3] = _zz_io_result_159[3];
    _zz_io_result_86[2] = _zz_io_result_159[2];
    _zz_io_result_86[1] = (! _zz_io_result_159[1]);
    _zz_io_result_86[0] = (! _zz_io_result_159[0]);
  end

  assign _zz_io_result_161 = _zz_io_result[23 : 16];
  always @(*) begin
    _zz_io_result_164[7] = (((((_zz_io_result_161[7] ^ _zz_io_result_161[6]) ^ _zz_io_result_161[5]) ^ _zz_io_result_161[2]) ^ _zz_io_result_161[1]) ^ _zz_io_result_161[0]);
    _zz_io_result_164[6] = (((_zz_io_result_161[6] ^ _zz_io_result_161[5]) ^ _zz_io_result_161[4]) ^ _zz_io_result_161[0]);
    _zz_io_result_164[5] = (((_zz_io_result_161[6] ^ _zz_io_result_161[5]) ^ _zz_io_result_161[1]) ^ _zz_io_result_161[0]);
    _zz_io_result_164[4] = (((_zz_io_result_161[7] ^ _zz_io_result_161[6]) ^ _zz_io_result_161[5]) ^ _zz_io_result_161[0]);
    _zz_io_result_164[3] = ((((_zz_io_result_161[7] ^ _zz_io_result_161[4]) ^ _zz_io_result_161[3]) ^ _zz_io_result_161[1]) ^ _zz_io_result_161[0]);
    _zz_io_result_164[2] = _zz_io_result_161[0];
    _zz_io_result_164[1] = ((_zz_io_result_161[6] ^ _zz_io_result_161[5]) ^ _zz_io_result_161[0]);
    _zz_io_result_164[0] = ((((_zz_io_result_161[6] ^ _zz_io_result_161[3]) ^ _zz_io_result_161[2]) ^ _zz_io_result_161[1]) ^ _zz_io_result_161[0]);
  end

  assign _zz_io_result_163 = _zz_io_result_164;
  assign _zz_io_result_167 = _zz_io_result_163[7 : 4];
  assign _zz_io_result_168 = _zz_io_result_163[3 : 0];
  assign _zz_io_result_169 = (_zz_io_result_167 ^ _zz_io_result_168);
  always @(*) begin
    _zz_io_result_170[3] = (_zz_io_result_169[2] ^ _zz_io_result_169[0]);
    _zz_io_result_170[2] = (_zz_io_result_169[3] ^ _zz_io_result_169[1]);
    _zz_io_result_170[1] = (_zz_io_result_169[1] ^ _zz_io_result_169[0]);
    _zz_io_result_170[0] = _zz_io_result_169[0];
  end

  assign _zz_io_result_172 = _zz_io_result_167[3 : 2];
  assign _zz_io_result_173 = _zz_io_result_167[1 : 0];
  assign _zz_io_result_174 = _zz_io_result_168[3 : 2];
  assign _zz_io_result_175 = _zz_io_result_168[1 : 0];
  assign _zz_io_result_176 = (_zz_io_result_172 ^ _zz_io_result_173);
  assign _zz_io_result_177 = (_zz_io_result_174 ^ _zz_io_result_175);
  assign _zz_io_result_179 = ((_zz_io_result_177[0] && _zz_io_result_176[1]) ^ (_zz_io_result_176[0] && _zz_io_result_177[1]));
  always @(*) begin
    _zz_io_result_180[1] = ((_zz_io_result_177[0] && _zz_io_result_176[0]) ^ _zz_io_result_179);
    _zz_io_result_180[0] = ((_zz_io_result_177[1] && _zz_io_result_176[1]) ^ _zz_io_result_179);
  end

  assign _zz_io_result_178 = _zz_io_result_180;
  always @(*) begin
    _zz_io_result_182[1] = _zz_io_result_178[0];
    _zz_io_result_182[0] = (_zz_io_result_178[0] ^ _zz_io_result_178[1]);
  end

  assign _zz_io_result_181 = _zz_io_result_182;
  assign _zz_io_result_183 = ((_zz_io_result_174[0] && _zz_io_result_172[1]) ^ (_zz_io_result_172[0] && _zz_io_result_174[1]));
  always @(*) begin
    _zz_io_result_184[1] = ((_zz_io_result_174[0] && _zz_io_result_172[0]) ^ _zz_io_result_183);
    _zz_io_result_184[0] = ((_zz_io_result_174[1] && _zz_io_result_172[1]) ^ _zz_io_result_183);
  end

  assign _zz_io_result_185 = ((_zz_io_result_175[0] && _zz_io_result_173[1]) ^ (_zz_io_result_173[0] && _zz_io_result_175[1]));
  always @(*) begin
    _zz_io_result_186[1] = ((_zz_io_result_175[0] && _zz_io_result_173[0]) ^ _zz_io_result_185);
    _zz_io_result_186[0] = ((_zz_io_result_175[1] && _zz_io_result_173[1]) ^ _zz_io_result_185);
  end

  always @(*) begin
    _zz_io_result_171[3 : 2] = (_zz_io_result_184 ^ _zz_io_result_181);
    _zz_io_result_171[1 : 0] = (_zz_io_result_186 ^ _zz_io_result_181);
  end

  assign _zz_io_result_187 = (_zz_io_result_170 ^ _zz_io_result_171);
  assign _zz_io_result_190 = _zz_io_result_187[3 : 2];
  assign _zz_io_result_191 = _zz_io_result_187[1 : 0];
  assign _zz_io_result_192 = (_zz_io_result_190 ^ _zz_io_result_191);
  always @(*) begin
    _zz_io_result_193[1] = _zz_io_result_192[1];
    _zz_io_result_193[0] = (_zz_io_result_192[0] ^ _zz_io_result_192[1]);
  end

  assign _zz_io_result_194 = ((_zz_io_result_191[0] && _zz_io_result_190[1]) ^ (_zz_io_result_190[0] && _zz_io_result_191[1]));
  always @(*) begin
    _zz_io_result_195[1] = ((_zz_io_result_191[0] && _zz_io_result_190[0]) ^ _zz_io_result_194);
    _zz_io_result_195[0] = ((_zz_io_result_191[1] && _zz_io_result_190[1]) ^ _zz_io_result_194);
  end

  assign _zz_io_result_196 = (_zz_io_result_193 ^ _zz_io_result_195);
  always @(*) begin
    _zz_io_result_198[1] = _zz_io_result_196[0];
    _zz_io_result_198[0] = _zz_io_result_196[1];
  end

  assign _zz_io_result_197 = _zz_io_result_198;
  assign _zz_io_result_199 = ((_zz_io_result_197[0] && _zz_io_result_190[1]) ^ (_zz_io_result_190[0] && _zz_io_result_197[1]));
  always @(*) begin
    _zz_io_result_200[1] = ((_zz_io_result_197[0] && _zz_io_result_190[0]) ^ _zz_io_result_199);
    _zz_io_result_200[0] = ((_zz_io_result_197[1] && _zz_io_result_190[1]) ^ _zz_io_result_199);
  end

  assign _zz_io_result_201 = ((_zz_io_result_197[0] && _zz_io_result_191[1]) ^ (_zz_io_result_191[0] && _zz_io_result_197[1]));
  always @(*) begin
    _zz_io_result_202[1] = ((_zz_io_result_197[0] && _zz_io_result_191[0]) ^ _zz_io_result_201);
    _zz_io_result_202[0] = ((_zz_io_result_197[1] && _zz_io_result_191[1]) ^ _zz_io_result_201);
  end

  always @(*) begin
    _zz_io_result_189[3 : 2] = _zz_io_result_202;
    _zz_io_result_189[1 : 0] = _zz_io_result_200;
  end

  assign _zz_io_result_188 = _zz_io_result_189;
  assign _zz_io_result_204 = _zz_io_result_167[3 : 2];
  assign _zz_io_result_205 = _zz_io_result_167[1 : 0];
  assign _zz_io_result_206 = _zz_io_result_188[3 : 2];
  assign _zz_io_result_207 = _zz_io_result_188[1 : 0];
  assign _zz_io_result_208 = (_zz_io_result_204 ^ _zz_io_result_205);
  assign _zz_io_result_209 = (_zz_io_result_206 ^ _zz_io_result_207);
  assign _zz_io_result_211 = ((_zz_io_result_209[0] && _zz_io_result_208[1]) ^ (_zz_io_result_208[0] && _zz_io_result_209[1]));
  always @(*) begin
    _zz_io_result_212[1] = ((_zz_io_result_209[0] && _zz_io_result_208[0]) ^ _zz_io_result_211);
    _zz_io_result_212[0] = ((_zz_io_result_209[1] && _zz_io_result_208[1]) ^ _zz_io_result_211);
  end

  assign _zz_io_result_210 = _zz_io_result_212;
  always @(*) begin
    _zz_io_result_214[1] = _zz_io_result_210[0];
    _zz_io_result_214[0] = (_zz_io_result_210[0] ^ _zz_io_result_210[1]);
  end

  assign _zz_io_result_213 = _zz_io_result_214;
  assign _zz_io_result_215 = ((_zz_io_result_206[0] && _zz_io_result_204[1]) ^ (_zz_io_result_204[0] && _zz_io_result_206[1]));
  always @(*) begin
    _zz_io_result_216[1] = ((_zz_io_result_206[0] && _zz_io_result_204[0]) ^ _zz_io_result_215);
    _zz_io_result_216[0] = ((_zz_io_result_206[1] && _zz_io_result_204[1]) ^ _zz_io_result_215);
  end

  assign _zz_io_result_217 = ((_zz_io_result_207[0] && _zz_io_result_205[1]) ^ (_zz_io_result_205[0] && _zz_io_result_207[1]));
  always @(*) begin
    _zz_io_result_218[1] = ((_zz_io_result_207[0] && _zz_io_result_205[0]) ^ _zz_io_result_217);
    _zz_io_result_218[0] = ((_zz_io_result_207[1] && _zz_io_result_205[1]) ^ _zz_io_result_217);
  end

  always @(*) begin
    _zz_io_result_203[3 : 2] = (_zz_io_result_216 ^ _zz_io_result_213);
    _zz_io_result_203[1 : 0] = (_zz_io_result_218 ^ _zz_io_result_213);
  end

  assign _zz_io_result_220 = _zz_io_result_168[3 : 2];
  assign _zz_io_result_221 = _zz_io_result_168[1 : 0];
  assign _zz_io_result_222 = _zz_io_result_188[3 : 2];
  assign _zz_io_result_223 = _zz_io_result_188[1 : 0];
  assign _zz_io_result_224 = (_zz_io_result_220 ^ _zz_io_result_221);
  assign _zz_io_result_225 = (_zz_io_result_222 ^ _zz_io_result_223);
  assign _zz_io_result_227 = ((_zz_io_result_225[0] && _zz_io_result_224[1]) ^ (_zz_io_result_224[0] && _zz_io_result_225[1]));
  always @(*) begin
    _zz_io_result_228[1] = ((_zz_io_result_225[0] && _zz_io_result_224[0]) ^ _zz_io_result_227);
    _zz_io_result_228[0] = ((_zz_io_result_225[1] && _zz_io_result_224[1]) ^ _zz_io_result_227);
  end

  assign _zz_io_result_226 = _zz_io_result_228;
  always @(*) begin
    _zz_io_result_230[1] = _zz_io_result_226[0];
    _zz_io_result_230[0] = (_zz_io_result_226[0] ^ _zz_io_result_226[1]);
  end

  assign _zz_io_result_229 = _zz_io_result_230;
  assign _zz_io_result_231 = ((_zz_io_result_222[0] && _zz_io_result_220[1]) ^ (_zz_io_result_220[0] && _zz_io_result_222[1]));
  always @(*) begin
    _zz_io_result_232[1] = ((_zz_io_result_222[0] && _zz_io_result_220[0]) ^ _zz_io_result_231);
    _zz_io_result_232[0] = ((_zz_io_result_222[1] && _zz_io_result_220[1]) ^ _zz_io_result_231);
  end

  assign _zz_io_result_233 = ((_zz_io_result_223[0] && _zz_io_result_221[1]) ^ (_zz_io_result_221[0] && _zz_io_result_223[1]));
  always @(*) begin
    _zz_io_result_234[1] = ((_zz_io_result_223[0] && _zz_io_result_221[0]) ^ _zz_io_result_233);
    _zz_io_result_234[0] = ((_zz_io_result_223[1] && _zz_io_result_221[1]) ^ _zz_io_result_233);
  end

  always @(*) begin
    _zz_io_result_219[3 : 2] = (_zz_io_result_232 ^ _zz_io_result_229);
    _zz_io_result_219[1 : 0] = (_zz_io_result_234 ^ _zz_io_result_229);
  end

  always @(*) begin
    _zz_io_result_166[7 : 4] = _zz_io_result_219;
    _zz_io_result_166[3 : 0] = _zz_io_result_203;
  end

  assign _zz_io_result_165 = _zz_io_result_166;
  always @(*) begin
    _zz_io_result_236[7] = (_zz_io_result_165[5] ^ _zz_io_result_165[3]);
    _zz_io_result_236[6] = (_zz_io_result_165[7] ^ _zz_io_result_165[3]);
    _zz_io_result_236[5] = (_zz_io_result_165[6] ^ _zz_io_result_165[0]);
    _zz_io_result_236[4] = ((_zz_io_result_165[7] ^ _zz_io_result_165[5]) ^ _zz_io_result_165[3]);
    _zz_io_result_236[3] = ((((_zz_io_result_165[7] ^ _zz_io_result_165[6]) ^ _zz_io_result_165[5]) ^ _zz_io_result_165[4]) ^ _zz_io_result_165[3]);
    _zz_io_result_236[2] = ((((_zz_io_result_165[6] ^ _zz_io_result_165[5]) ^ _zz_io_result_165[3]) ^ _zz_io_result_165[2]) ^ _zz_io_result_165[0]);
    _zz_io_result_236[1] = ((_zz_io_result_165[5] ^ _zz_io_result_165[4]) ^ _zz_io_result_165[1]);
    _zz_io_result_236[0] = ((_zz_io_result_165[6] ^ _zz_io_result_165[4]) ^ _zz_io_result_165[1]);
  end

  assign _zz_io_result_235 = _zz_io_result_236;
  always @(*) begin
    _zz_io_result_162[7] = _zz_io_result_235[7];
    _zz_io_result_162[6] = (! _zz_io_result_235[6]);
    _zz_io_result_162[5] = (! _zz_io_result_235[5]);
    _zz_io_result_162[4] = _zz_io_result_235[4];
    _zz_io_result_162[3] = _zz_io_result_235[3];
    _zz_io_result_162[2] = _zz_io_result_235[2];
    _zz_io_result_162[1] = (! _zz_io_result_235[1]);
    _zz_io_result_162[0] = (! _zz_io_result_235[0]);
  end

  assign _zz_io_result_237 = _zz_io_result[31 : 24];
  always @(*) begin
    _zz_io_result_240[7] = (((((_zz_io_result_237[7] ^ _zz_io_result_237[6]) ^ _zz_io_result_237[5]) ^ _zz_io_result_237[2]) ^ _zz_io_result_237[1]) ^ _zz_io_result_237[0]);
    _zz_io_result_240[6] = (((_zz_io_result_237[6] ^ _zz_io_result_237[5]) ^ _zz_io_result_237[4]) ^ _zz_io_result_237[0]);
    _zz_io_result_240[5] = (((_zz_io_result_237[6] ^ _zz_io_result_237[5]) ^ _zz_io_result_237[1]) ^ _zz_io_result_237[0]);
    _zz_io_result_240[4] = (((_zz_io_result_237[7] ^ _zz_io_result_237[6]) ^ _zz_io_result_237[5]) ^ _zz_io_result_237[0]);
    _zz_io_result_240[3] = ((((_zz_io_result_237[7] ^ _zz_io_result_237[4]) ^ _zz_io_result_237[3]) ^ _zz_io_result_237[1]) ^ _zz_io_result_237[0]);
    _zz_io_result_240[2] = _zz_io_result_237[0];
    _zz_io_result_240[1] = ((_zz_io_result_237[6] ^ _zz_io_result_237[5]) ^ _zz_io_result_237[0]);
    _zz_io_result_240[0] = ((((_zz_io_result_237[6] ^ _zz_io_result_237[3]) ^ _zz_io_result_237[2]) ^ _zz_io_result_237[1]) ^ _zz_io_result_237[0]);
  end

  assign _zz_io_result_239 = _zz_io_result_240;
  assign _zz_io_result_243 = _zz_io_result_239[7 : 4];
  assign _zz_io_result_244 = _zz_io_result_239[3 : 0];
  assign _zz_io_result_245 = (_zz_io_result_243 ^ _zz_io_result_244);
  always @(*) begin
    _zz_io_result_246[3] = (_zz_io_result_245[2] ^ _zz_io_result_245[0]);
    _zz_io_result_246[2] = (_zz_io_result_245[3] ^ _zz_io_result_245[1]);
    _zz_io_result_246[1] = (_zz_io_result_245[1] ^ _zz_io_result_245[0]);
    _zz_io_result_246[0] = _zz_io_result_245[0];
  end

  assign _zz_io_result_248 = _zz_io_result_243[3 : 2];
  assign _zz_io_result_249 = _zz_io_result_243[1 : 0];
  assign _zz_io_result_250 = _zz_io_result_244[3 : 2];
  assign _zz_io_result_251 = _zz_io_result_244[1 : 0];
  assign _zz_io_result_252 = (_zz_io_result_248 ^ _zz_io_result_249);
  assign _zz_io_result_253 = (_zz_io_result_250 ^ _zz_io_result_251);
  assign _zz_io_result_255 = ((_zz_io_result_253[0] && _zz_io_result_252[1]) ^ (_zz_io_result_252[0] && _zz_io_result_253[1]));
  always @(*) begin
    _zz_io_result_256[1] = ((_zz_io_result_253[0] && _zz_io_result_252[0]) ^ _zz_io_result_255);
    _zz_io_result_256[0] = ((_zz_io_result_253[1] && _zz_io_result_252[1]) ^ _zz_io_result_255);
  end

  assign _zz_io_result_254 = _zz_io_result_256;
  always @(*) begin
    _zz_io_result_258[1] = _zz_io_result_254[0];
    _zz_io_result_258[0] = (_zz_io_result_254[0] ^ _zz_io_result_254[1]);
  end

  assign _zz_io_result_257 = _zz_io_result_258;
  assign _zz_io_result_259 = ((_zz_io_result_250[0] && _zz_io_result_248[1]) ^ (_zz_io_result_248[0] && _zz_io_result_250[1]));
  always @(*) begin
    _zz_io_result_260[1] = ((_zz_io_result_250[0] && _zz_io_result_248[0]) ^ _zz_io_result_259);
    _zz_io_result_260[0] = ((_zz_io_result_250[1] && _zz_io_result_248[1]) ^ _zz_io_result_259);
  end

  assign _zz_io_result_261 = ((_zz_io_result_251[0] && _zz_io_result_249[1]) ^ (_zz_io_result_249[0] && _zz_io_result_251[1]));
  always @(*) begin
    _zz_io_result_262[1] = ((_zz_io_result_251[0] && _zz_io_result_249[0]) ^ _zz_io_result_261);
    _zz_io_result_262[0] = ((_zz_io_result_251[1] && _zz_io_result_249[1]) ^ _zz_io_result_261);
  end

  always @(*) begin
    _zz_io_result_247[3 : 2] = (_zz_io_result_260 ^ _zz_io_result_257);
    _zz_io_result_247[1 : 0] = (_zz_io_result_262 ^ _zz_io_result_257);
  end

  assign _zz_io_result_263 = (_zz_io_result_246 ^ _zz_io_result_247);
  assign _zz_io_result_266 = _zz_io_result_263[3 : 2];
  assign _zz_io_result_267 = _zz_io_result_263[1 : 0];
  assign _zz_io_result_268 = (_zz_io_result_266 ^ _zz_io_result_267);
  always @(*) begin
    _zz_io_result_269[1] = _zz_io_result_268[1];
    _zz_io_result_269[0] = (_zz_io_result_268[0] ^ _zz_io_result_268[1]);
  end

  assign _zz_io_result_270 = ((_zz_io_result_267[0] && _zz_io_result_266[1]) ^ (_zz_io_result_266[0] && _zz_io_result_267[1]));
  always @(*) begin
    _zz_io_result_271[1] = ((_zz_io_result_267[0] && _zz_io_result_266[0]) ^ _zz_io_result_270);
    _zz_io_result_271[0] = ((_zz_io_result_267[1] && _zz_io_result_266[1]) ^ _zz_io_result_270);
  end

  assign _zz_io_result_272 = (_zz_io_result_269 ^ _zz_io_result_271);
  always @(*) begin
    _zz_io_result_274[1] = _zz_io_result_272[0];
    _zz_io_result_274[0] = _zz_io_result_272[1];
  end

  assign _zz_io_result_273 = _zz_io_result_274;
  assign _zz_io_result_275 = ((_zz_io_result_273[0] && _zz_io_result_266[1]) ^ (_zz_io_result_266[0] && _zz_io_result_273[1]));
  always @(*) begin
    _zz_io_result_276[1] = ((_zz_io_result_273[0] && _zz_io_result_266[0]) ^ _zz_io_result_275);
    _zz_io_result_276[0] = ((_zz_io_result_273[1] && _zz_io_result_266[1]) ^ _zz_io_result_275);
  end

  assign _zz_io_result_277 = ((_zz_io_result_273[0] && _zz_io_result_267[1]) ^ (_zz_io_result_267[0] && _zz_io_result_273[1]));
  always @(*) begin
    _zz_io_result_278[1] = ((_zz_io_result_273[0] && _zz_io_result_267[0]) ^ _zz_io_result_277);
    _zz_io_result_278[0] = ((_zz_io_result_273[1] && _zz_io_result_267[1]) ^ _zz_io_result_277);
  end

  always @(*) begin
    _zz_io_result_265[3 : 2] = _zz_io_result_278;
    _zz_io_result_265[1 : 0] = _zz_io_result_276;
  end

  assign _zz_io_result_264 = _zz_io_result_265;
  assign _zz_io_result_280 = _zz_io_result_243[3 : 2];
  assign _zz_io_result_281 = _zz_io_result_243[1 : 0];
  assign _zz_io_result_282 = _zz_io_result_264[3 : 2];
  assign _zz_io_result_283 = _zz_io_result_264[1 : 0];
  assign _zz_io_result_284 = (_zz_io_result_280 ^ _zz_io_result_281);
  assign _zz_io_result_285 = (_zz_io_result_282 ^ _zz_io_result_283);
  assign _zz_io_result_287 = ((_zz_io_result_285[0] && _zz_io_result_284[1]) ^ (_zz_io_result_284[0] && _zz_io_result_285[1]));
  always @(*) begin
    _zz_io_result_288[1] = ((_zz_io_result_285[0] && _zz_io_result_284[0]) ^ _zz_io_result_287);
    _zz_io_result_288[0] = ((_zz_io_result_285[1] && _zz_io_result_284[1]) ^ _zz_io_result_287);
  end

  assign _zz_io_result_286 = _zz_io_result_288;
  always @(*) begin
    _zz_io_result_290[1] = _zz_io_result_286[0];
    _zz_io_result_290[0] = (_zz_io_result_286[0] ^ _zz_io_result_286[1]);
  end

  assign _zz_io_result_289 = _zz_io_result_290;
  assign _zz_io_result_291 = ((_zz_io_result_282[0] && _zz_io_result_280[1]) ^ (_zz_io_result_280[0] && _zz_io_result_282[1]));
  always @(*) begin
    _zz_io_result_292[1] = ((_zz_io_result_282[0] && _zz_io_result_280[0]) ^ _zz_io_result_291);
    _zz_io_result_292[0] = ((_zz_io_result_282[1] && _zz_io_result_280[1]) ^ _zz_io_result_291);
  end

  assign _zz_io_result_293 = ((_zz_io_result_283[0] && _zz_io_result_281[1]) ^ (_zz_io_result_281[0] && _zz_io_result_283[1]));
  always @(*) begin
    _zz_io_result_294[1] = ((_zz_io_result_283[0] && _zz_io_result_281[0]) ^ _zz_io_result_293);
    _zz_io_result_294[0] = ((_zz_io_result_283[1] && _zz_io_result_281[1]) ^ _zz_io_result_293);
  end

  always @(*) begin
    _zz_io_result_279[3 : 2] = (_zz_io_result_292 ^ _zz_io_result_289);
    _zz_io_result_279[1 : 0] = (_zz_io_result_294 ^ _zz_io_result_289);
  end

  assign _zz_io_result_296 = _zz_io_result_244[3 : 2];
  assign _zz_io_result_297 = _zz_io_result_244[1 : 0];
  assign _zz_io_result_298 = _zz_io_result_264[3 : 2];
  assign _zz_io_result_299 = _zz_io_result_264[1 : 0];
  assign _zz_io_result_300 = (_zz_io_result_296 ^ _zz_io_result_297);
  assign _zz_io_result_301 = (_zz_io_result_298 ^ _zz_io_result_299);
  assign _zz_io_result_303 = ((_zz_io_result_301[0] && _zz_io_result_300[1]) ^ (_zz_io_result_300[0] && _zz_io_result_301[1]));
  always @(*) begin
    _zz_io_result_304[1] = ((_zz_io_result_301[0] && _zz_io_result_300[0]) ^ _zz_io_result_303);
    _zz_io_result_304[0] = ((_zz_io_result_301[1] && _zz_io_result_300[1]) ^ _zz_io_result_303);
  end

  assign _zz_io_result_302 = _zz_io_result_304;
  always @(*) begin
    _zz_io_result_306[1] = _zz_io_result_302[0];
    _zz_io_result_306[0] = (_zz_io_result_302[0] ^ _zz_io_result_302[1]);
  end

  assign _zz_io_result_305 = _zz_io_result_306;
  assign _zz_io_result_307 = ((_zz_io_result_298[0] && _zz_io_result_296[1]) ^ (_zz_io_result_296[0] && _zz_io_result_298[1]));
  always @(*) begin
    _zz_io_result_308[1] = ((_zz_io_result_298[0] && _zz_io_result_296[0]) ^ _zz_io_result_307);
    _zz_io_result_308[0] = ((_zz_io_result_298[1] && _zz_io_result_296[1]) ^ _zz_io_result_307);
  end

  assign _zz_io_result_309 = ((_zz_io_result_299[0] && _zz_io_result_297[1]) ^ (_zz_io_result_297[0] && _zz_io_result_299[1]));
  always @(*) begin
    _zz_io_result_310[1] = ((_zz_io_result_299[0] && _zz_io_result_297[0]) ^ _zz_io_result_309);
    _zz_io_result_310[0] = ((_zz_io_result_299[1] && _zz_io_result_297[1]) ^ _zz_io_result_309);
  end

  always @(*) begin
    _zz_io_result_295[3 : 2] = (_zz_io_result_308 ^ _zz_io_result_305);
    _zz_io_result_295[1 : 0] = (_zz_io_result_310 ^ _zz_io_result_305);
  end

  always @(*) begin
    _zz_io_result_242[7 : 4] = _zz_io_result_295;
    _zz_io_result_242[3 : 0] = _zz_io_result_279;
  end

  assign _zz_io_result_241 = _zz_io_result_242;
  always @(*) begin
    _zz_io_result_312[7] = (_zz_io_result_241[5] ^ _zz_io_result_241[3]);
    _zz_io_result_312[6] = (_zz_io_result_241[7] ^ _zz_io_result_241[3]);
    _zz_io_result_312[5] = (_zz_io_result_241[6] ^ _zz_io_result_241[0]);
    _zz_io_result_312[4] = ((_zz_io_result_241[7] ^ _zz_io_result_241[5]) ^ _zz_io_result_241[3]);
    _zz_io_result_312[3] = ((((_zz_io_result_241[7] ^ _zz_io_result_241[6]) ^ _zz_io_result_241[5]) ^ _zz_io_result_241[4]) ^ _zz_io_result_241[3]);
    _zz_io_result_312[2] = ((((_zz_io_result_241[6] ^ _zz_io_result_241[5]) ^ _zz_io_result_241[3]) ^ _zz_io_result_241[2]) ^ _zz_io_result_241[0]);
    _zz_io_result_312[1] = ((_zz_io_result_241[5] ^ _zz_io_result_241[4]) ^ _zz_io_result_241[1]);
    _zz_io_result_312[0] = ((_zz_io_result_241[6] ^ _zz_io_result_241[4]) ^ _zz_io_result_241[1]);
  end

  assign _zz_io_result_311 = _zz_io_result_312;
  always @(*) begin
    _zz_io_result_238[7] = _zz_io_result_311[7];
    _zz_io_result_238[6] = (! _zz_io_result_311[6]);
    _zz_io_result_238[5] = (! _zz_io_result_311[5]);
    _zz_io_result_238[4] = _zz_io_result_311[4];
    _zz_io_result_238[3] = _zz_io_result_311[3];
    _zz_io_result_238[2] = _zz_io_result_311[2];
    _zz_io_result_238[1] = (! _zz_io_result_311[1]);
    _zz_io_result_238[0] = (! _zz_io_result_311[0]);
  end

  assign _zz_io_result_314 = _zz_io_result_1[7 : 0];
  always @(*) begin
    _zz_io_result_317[7] = (((((_zz_io_result_314[7] ^ _zz_io_result_314[6]) ^ _zz_io_result_314[5]) ^ _zz_io_result_314[2]) ^ _zz_io_result_314[1]) ^ _zz_io_result_314[0]);
    _zz_io_result_317[6] = (((_zz_io_result_314[6] ^ _zz_io_result_314[5]) ^ _zz_io_result_314[4]) ^ _zz_io_result_314[0]);
    _zz_io_result_317[5] = (((_zz_io_result_314[6] ^ _zz_io_result_314[5]) ^ _zz_io_result_314[1]) ^ _zz_io_result_314[0]);
    _zz_io_result_317[4] = (((_zz_io_result_314[7] ^ _zz_io_result_314[6]) ^ _zz_io_result_314[5]) ^ _zz_io_result_314[0]);
    _zz_io_result_317[3] = ((((_zz_io_result_314[7] ^ _zz_io_result_314[4]) ^ _zz_io_result_314[3]) ^ _zz_io_result_314[1]) ^ _zz_io_result_314[0]);
    _zz_io_result_317[2] = _zz_io_result_314[0];
    _zz_io_result_317[1] = ((_zz_io_result_314[6] ^ _zz_io_result_314[5]) ^ _zz_io_result_314[0]);
    _zz_io_result_317[0] = ((((_zz_io_result_314[6] ^ _zz_io_result_314[3]) ^ _zz_io_result_314[2]) ^ _zz_io_result_314[1]) ^ _zz_io_result_314[0]);
  end

  assign _zz_io_result_316 = _zz_io_result_317;
  assign _zz_io_result_320 = _zz_io_result_316[7 : 4];
  assign _zz_io_result_321 = _zz_io_result_316[3 : 0];
  assign _zz_io_result_322 = (_zz_io_result_320 ^ _zz_io_result_321);
  always @(*) begin
    _zz_io_result_323[3] = (_zz_io_result_322[2] ^ _zz_io_result_322[0]);
    _zz_io_result_323[2] = (_zz_io_result_322[3] ^ _zz_io_result_322[1]);
    _zz_io_result_323[1] = (_zz_io_result_322[1] ^ _zz_io_result_322[0]);
    _zz_io_result_323[0] = _zz_io_result_322[0];
  end

  assign _zz_io_result_325 = _zz_io_result_320[3 : 2];
  assign _zz_io_result_326 = _zz_io_result_320[1 : 0];
  assign _zz_io_result_327 = _zz_io_result_321[3 : 2];
  assign _zz_io_result_328 = _zz_io_result_321[1 : 0];
  assign _zz_io_result_329 = (_zz_io_result_325 ^ _zz_io_result_326);
  assign _zz_io_result_330 = (_zz_io_result_327 ^ _zz_io_result_328);
  assign _zz_io_result_332 = ((_zz_io_result_330[0] && _zz_io_result_329[1]) ^ (_zz_io_result_329[0] && _zz_io_result_330[1]));
  always @(*) begin
    _zz_io_result_333[1] = ((_zz_io_result_330[0] && _zz_io_result_329[0]) ^ _zz_io_result_332);
    _zz_io_result_333[0] = ((_zz_io_result_330[1] && _zz_io_result_329[1]) ^ _zz_io_result_332);
  end

  assign _zz_io_result_331 = _zz_io_result_333;
  always @(*) begin
    _zz_io_result_335[1] = _zz_io_result_331[0];
    _zz_io_result_335[0] = (_zz_io_result_331[0] ^ _zz_io_result_331[1]);
  end

  assign _zz_io_result_334 = _zz_io_result_335;
  assign _zz_io_result_336 = ((_zz_io_result_327[0] && _zz_io_result_325[1]) ^ (_zz_io_result_325[0] && _zz_io_result_327[1]));
  always @(*) begin
    _zz_io_result_337[1] = ((_zz_io_result_327[0] && _zz_io_result_325[0]) ^ _zz_io_result_336);
    _zz_io_result_337[0] = ((_zz_io_result_327[1] && _zz_io_result_325[1]) ^ _zz_io_result_336);
  end

  assign _zz_io_result_338 = ((_zz_io_result_328[0] && _zz_io_result_326[1]) ^ (_zz_io_result_326[0] && _zz_io_result_328[1]));
  always @(*) begin
    _zz_io_result_339[1] = ((_zz_io_result_328[0] && _zz_io_result_326[0]) ^ _zz_io_result_338);
    _zz_io_result_339[0] = ((_zz_io_result_328[1] && _zz_io_result_326[1]) ^ _zz_io_result_338);
  end

  always @(*) begin
    _zz_io_result_324[3 : 2] = (_zz_io_result_337 ^ _zz_io_result_334);
    _zz_io_result_324[1 : 0] = (_zz_io_result_339 ^ _zz_io_result_334);
  end

  assign _zz_io_result_340 = (_zz_io_result_323 ^ _zz_io_result_324);
  assign _zz_io_result_343 = _zz_io_result_340[3 : 2];
  assign _zz_io_result_344 = _zz_io_result_340[1 : 0];
  assign _zz_io_result_345 = (_zz_io_result_343 ^ _zz_io_result_344);
  always @(*) begin
    _zz_io_result_346[1] = _zz_io_result_345[1];
    _zz_io_result_346[0] = (_zz_io_result_345[0] ^ _zz_io_result_345[1]);
  end

  assign _zz_io_result_347 = ((_zz_io_result_344[0] && _zz_io_result_343[1]) ^ (_zz_io_result_343[0] && _zz_io_result_344[1]));
  always @(*) begin
    _zz_io_result_348[1] = ((_zz_io_result_344[0] && _zz_io_result_343[0]) ^ _zz_io_result_347);
    _zz_io_result_348[0] = ((_zz_io_result_344[1] && _zz_io_result_343[1]) ^ _zz_io_result_347);
  end

  assign _zz_io_result_349 = (_zz_io_result_346 ^ _zz_io_result_348);
  always @(*) begin
    _zz_io_result_351[1] = _zz_io_result_349[0];
    _zz_io_result_351[0] = _zz_io_result_349[1];
  end

  assign _zz_io_result_350 = _zz_io_result_351;
  assign _zz_io_result_352 = ((_zz_io_result_350[0] && _zz_io_result_343[1]) ^ (_zz_io_result_343[0] && _zz_io_result_350[1]));
  always @(*) begin
    _zz_io_result_353[1] = ((_zz_io_result_350[0] && _zz_io_result_343[0]) ^ _zz_io_result_352);
    _zz_io_result_353[0] = ((_zz_io_result_350[1] && _zz_io_result_343[1]) ^ _zz_io_result_352);
  end

  assign _zz_io_result_354 = ((_zz_io_result_350[0] && _zz_io_result_344[1]) ^ (_zz_io_result_344[0] && _zz_io_result_350[1]));
  always @(*) begin
    _zz_io_result_355[1] = ((_zz_io_result_350[0] && _zz_io_result_344[0]) ^ _zz_io_result_354);
    _zz_io_result_355[0] = ((_zz_io_result_350[1] && _zz_io_result_344[1]) ^ _zz_io_result_354);
  end

  always @(*) begin
    _zz_io_result_342[3 : 2] = _zz_io_result_355;
    _zz_io_result_342[1 : 0] = _zz_io_result_353;
  end

  assign _zz_io_result_341 = _zz_io_result_342;
  assign _zz_io_result_357 = _zz_io_result_320[3 : 2];
  assign _zz_io_result_358 = _zz_io_result_320[1 : 0];
  assign _zz_io_result_359 = _zz_io_result_341[3 : 2];
  assign _zz_io_result_360 = _zz_io_result_341[1 : 0];
  assign _zz_io_result_361 = (_zz_io_result_357 ^ _zz_io_result_358);
  assign _zz_io_result_362 = (_zz_io_result_359 ^ _zz_io_result_360);
  assign _zz_io_result_364 = ((_zz_io_result_362[0] && _zz_io_result_361[1]) ^ (_zz_io_result_361[0] && _zz_io_result_362[1]));
  always @(*) begin
    _zz_io_result_365[1] = ((_zz_io_result_362[0] && _zz_io_result_361[0]) ^ _zz_io_result_364);
    _zz_io_result_365[0] = ((_zz_io_result_362[1] && _zz_io_result_361[1]) ^ _zz_io_result_364);
  end

  assign _zz_io_result_363 = _zz_io_result_365;
  always @(*) begin
    _zz_io_result_367[1] = _zz_io_result_363[0];
    _zz_io_result_367[0] = (_zz_io_result_363[0] ^ _zz_io_result_363[1]);
  end

  assign _zz_io_result_366 = _zz_io_result_367;
  assign _zz_io_result_368 = ((_zz_io_result_359[0] && _zz_io_result_357[1]) ^ (_zz_io_result_357[0] && _zz_io_result_359[1]));
  always @(*) begin
    _zz_io_result_369[1] = ((_zz_io_result_359[0] && _zz_io_result_357[0]) ^ _zz_io_result_368);
    _zz_io_result_369[0] = ((_zz_io_result_359[1] && _zz_io_result_357[1]) ^ _zz_io_result_368);
  end

  assign _zz_io_result_370 = ((_zz_io_result_360[0] && _zz_io_result_358[1]) ^ (_zz_io_result_358[0] && _zz_io_result_360[1]));
  always @(*) begin
    _zz_io_result_371[1] = ((_zz_io_result_360[0] && _zz_io_result_358[0]) ^ _zz_io_result_370);
    _zz_io_result_371[0] = ((_zz_io_result_360[1] && _zz_io_result_358[1]) ^ _zz_io_result_370);
  end

  always @(*) begin
    _zz_io_result_356[3 : 2] = (_zz_io_result_369 ^ _zz_io_result_366);
    _zz_io_result_356[1 : 0] = (_zz_io_result_371 ^ _zz_io_result_366);
  end

  assign _zz_io_result_373 = _zz_io_result_321[3 : 2];
  assign _zz_io_result_374 = _zz_io_result_321[1 : 0];
  assign _zz_io_result_375 = _zz_io_result_341[3 : 2];
  assign _zz_io_result_376 = _zz_io_result_341[1 : 0];
  assign _zz_io_result_377 = (_zz_io_result_373 ^ _zz_io_result_374);
  assign _zz_io_result_378 = (_zz_io_result_375 ^ _zz_io_result_376);
  assign _zz_io_result_380 = ((_zz_io_result_378[0] && _zz_io_result_377[1]) ^ (_zz_io_result_377[0] && _zz_io_result_378[1]));
  always @(*) begin
    _zz_io_result_381[1] = ((_zz_io_result_378[0] && _zz_io_result_377[0]) ^ _zz_io_result_380);
    _zz_io_result_381[0] = ((_zz_io_result_378[1] && _zz_io_result_377[1]) ^ _zz_io_result_380);
  end

  assign _zz_io_result_379 = _zz_io_result_381;
  always @(*) begin
    _zz_io_result_383[1] = _zz_io_result_379[0];
    _zz_io_result_383[0] = (_zz_io_result_379[0] ^ _zz_io_result_379[1]);
  end

  assign _zz_io_result_382 = _zz_io_result_383;
  assign _zz_io_result_384 = ((_zz_io_result_375[0] && _zz_io_result_373[1]) ^ (_zz_io_result_373[0] && _zz_io_result_375[1]));
  always @(*) begin
    _zz_io_result_385[1] = ((_zz_io_result_375[0] && _zz_io_result_373[0]) ^ _zz_io_result_384);
    _zz_io_result_385[0] = ((_zz_io_result_375[1] && _zz_io_result_373[1]) ^ _zz_io_result_384);
  end

  assign _zz_io_result_386 = ((_zz_io_result_376[0] && _zz_io_result_374[1]) ^ (_zz_io_result_374[0] && _zz_io_result_376[1]));
  always @(*) begin
    _zz_io_result_387[1] = ((_zz_io_result_376[0] && _zz_io_result_374[0]) ^ _zz_io_result_386);
    _zz_io_result_387[0] = ((_zz_io_result_376[1] && _zz_io_result_374[1]) ^ _zz_io_result_386);
  end

  always @(*) begin
    _zz_io_result_372[3 : 2] = (_zz_io_result_385 ^ _zz_io_result_382);
    _zz_io_result_372[1 : 0] = (_zz_io_result_387 ^ _zz_io_result_382);
  end

  always @(*) begin
    _zz_io_result_319[7 : 4] = _zz_io_result_372;
    _zz_io_result_319[3 : 0] = _zz_io_result_356;
  end

  assign _zz_io_result_318 = _zz_io_result_319;
  always @(*) begin
    _zz_io_result_389[7] = (_zz_io_result_318[5] ^ _zz_io_result_318[3]);
    _zz_io_result_389[6] = (_zz_io_result_318[7] ^ _zz_io_result_318[3]);
    _zz_io_result_389[5] = (_zz_io_result_318[6] ^ _zz_io_result_318[0]);
    _zz_io_result_389[4] = ((_zz_io_result_318[7] ^ _zz_io_result_318[5]) ^ _zz_io_result_318[3]);
    _zz_io_result_389[3] = ((((_zz_io_result_318[7] ^ _zz_io_result_318[6]) ^ _zz_io_result_318[5]) ^ _zz_io_result_318[4]) ^ _zz_io_result_318[3]);
    _zz_io_result_389[2] = ((((_zz_io_result_318[6] ^ _zz_io_result_318[5]) ^ _zz_io_result_318[3]) ^ _zz_io_result_318[2]) ^ _zz_io_result_318[0]);
    _zz_io_result_389[1] = ((_zz_io_result_318[5] ^ _zz_io_result_318[4]) ^ _zz_io_result_318[1]);
    _zz_io_result_389[0] = ((_zz_io_result_318[6] ^ _zz_io_result_318[4]) ^ _zz_io_result_318[1]);
  end

  assign _zz_io_result_388 = _zz_io_result_389;
  always @(*) begin
    _zz_io_result_315[7] = _zz_io_result_388[7];
    _zz_io_result_315[6] = (! _zz_io_result_388[6]);
    _zz_io_result_315[5] = (! _zz_io_result_388[5]);
    _zz_io_result_315[4] = _zz_io_result_388[4];
    _zz_io_result_315[3] = _zz_io_result_388[3];
    _zz_io_result_315[2] = _zz_io_result_388[2];
    _zz_io_result_315[1] = (! _zz_io_result_388[1]);
    _zz_io_result_315[0] = (! _zz_io_result_388[0]);
  end

  always @(*) begin
    _zz_io_result_313[7 : 0] = _zz_io_result_315;
    _zz_io_result_313[15 : 8] = _zz_io_result_391;
    _zz_io_result_313[23 : 16] = _zz_io_result_467;
    _zz_io_result_313[31 : 24] = _zz_io_result_543;
  end

  assign _zz_io_result_390 = _zz_io_result_1[15 : 8];
  always @(*) begin
    _zz_io_result_393[7] = (((((_zz_io_result_390[7] ^ _zz_io_result_390[6]) ^ _zz_io_result_390[5]) ^ _zz_io_result_390[2]) ^ _zz_io_result_390[1]) ^ _zz_io_result_390[0]);
    _zz_io_result_393[6] = (((_zz_io_result_390[6] ^ _zz_io_result_390[5]) ^ _zz_io_result_390[4]) ^ _zz_io_result_390[0]);
    _zz_io_result_393[5] = (((_zz_io_result_390[6] ^ _zz_io_result_390[5]) ^ _zz_io_result_390[1]) ^ _zz_io_result_390[0]);
    _zz_io_result_393[4] = (((_zz_io_result_390[7] ^ _zz_io_result_390[6]) ^ _zz_io_result_390[5]) ^ _zz_io_result_390[0]);
    _zz_io_result_393[3] = ((((_zz_io_result_390[7] ^ _zz_io_result_390[4]) ^ _zz_io_result_390[3]) ^ _zz_io_result_390[1]) ^ _zz_io_result_390[0]);
    _zz_io_result_393[2] = _zz_io_result_390[0];
    _zz_io_result_393[1] = ((_zz_io_result_390[6] ^ _zz_io_result_390[5]) ^ _zz_io_result_390[0]);
    _zz_io_result_393[0] = ((((_zz_io_result_390[6] ^ _zz_io_result_390[3]) ^ _zz_io_result_390[2]) ^ _zz_io_result_390[1]) ^ _zz_io_result_390[0]);
  end

  assign _zz_io_result_392 = _zz_io_result_393;
  assign _zz_io_result_396 = _zz_io_result_392[7 : 4];
  assign _zz_io_result_397 = _zz_io_result_392[3 : 0];
  assign _zz_io_result_398 = (_zz_io_result_396 ^ _zz_io_result_397);
  always @(*) begin
    _zz_io_result_399[3] = (_zz_io_result_398[2] ^ _zz_io_result_398[0]);
    _zz_io_result_399[2] = (_zz_io_result_398[3] ^ _zz_io_result_398[1]);
    _zz_io_result_399[1] = (_zz_io_result_398[1] ^ _zz_io_result_398[0]);
    _zz_io_result_399[0] = _zz_io_result_398[0];
  end

  assign _zz_io_result_401 = _zz_io_result_396[3 : 2];
  assign _zz_io_result_402 = _zz_io_result_396[1 : 0];
  assign _zz_io_result_403 = _zz_io_result_397[3 : 2];
  assign _zz_io_result_404 = _zz_io_result_397[1 : 0];
  assign _zz_io_result_405 = (_zz_io_result_401 ^ _zz_io_result_402);
  assign _zz_io_result_406 = (_zz_io_result_403 ^ _zz_io_result_404);
  assign _zz_io_result_408 = ((_zz_io_result_406[0] && _zz_io_result_405[1]) ^ (_zz_io_result_405[0] && _zz_io_result_406[1]));
  always @(*) begin
    _zz_io_result_409[1] = ((_zz_io_result_406[0] && _zz_io_result_405[0]) ^ _zz_io_result_408);
    _zz_io_result_409[0] = ((_zz_io_result_406[1] && _zz_io_result_405[1]) ^ _zz_io_result_408);
  end

  assign _zz_io_result_407 = _zz_io_result_409;
  always @(*) begin
    _zz_io_result_411[1] = _zz_io_result_407[0];
    _zz_io_result_411[0] = (_zz_io_result_407[0] ^ _zz_io_result_407[1]);
  end

  assign _zz_io_result_410 = _zz_io_result_411;
  assign _zz_io_result_412 = ((_zz_io_result_403[0] && _zz_io_result_401[1]) ^ (_zz_io_result_401[0] && _zz_io_result_403[1]));
  always @(*) begin
    _zz_io_result_413[1] = ((_zz_io_result_403[0] && _zz_io_result_401[0]) ^ _zz_io_result_412);
    _zz_io_result_413[0] = ((_zz_io_result_403[1] && _zz_io_result_401[1]) ^ _zz_io_result_412);
  end

  assign _zz_io_result_414 = ((_zz_io_result_404[0] && _zz_io_result_402[1]) ^ (_zz_io_result_402[0] && _zz_io_result_404[1]));
  always @(*) begin
    _zz_io_result_415[1] = ((_zz_io_result_404[0] && _zz_io_result_402[0]) ^ _zz_io_result_414);
    _zz_io_result_415[0] = ((_zz_io_result_404[1] && _zz_io_result_402[1]) ^ _zz_io_result_414);
  end

  always @(*) begin
    _zz_io_result_400[3 : 2] = (_zz_io_result_413 ^ _zz_io_result_410);
    _zz_io_result_400[1 : 0] = (_zz_io_result_415 ^ _zz_io_result_410);
  end

  assign _zz_io_result_416 = (_zz_io_result_399 ^ _zz_io_result_400);
  assign _zz_io_result_419 = _zz_io_result_416[3 : 2];
  assign _zz_io_result_420 = _zz_io_result_416[1 : 0];
  assign _zz_io_result_421 = (_zz_io_result_419 ^ _zz_io_result_420);
  always @(*) begin
    _zz_io_result_422[1] = _zz_io_result_421[1];
    _zz_io_result_422[0] = (_zz_io_result_421[0] ^ _zz_io_result_421[1]);
  end

  assign _zz_io_result_423 = ((_zz_io_result_420[0] && _zz_io_result_419[1]) ^ (_zz_io_result_419[0] && _zz_io_result_420[1]));
  always @(*) begin
    _zz_io_result_424[1] = ((_zz_io_result_420[0] && _zz_io_result_419[0]) ^ _zz_io_result_423);
    _zz_io_result_424[0] = ((_zz_io_result_420[1] && _zz_io_result_419[1]) ^ _zz_io_result_423);
  end

  assign _zz_io_result_425 = (_zz_io_result_422 ^ _zz_io_result_424);
  always @(*) begin
    _zz_io_result_427[1] = _zz_io_result_425[0];
    _zz_io_result_427[0] = _zz_io_result_425[1];
  end

  assign _zz_io_result_426 = _zz_io_result_427;
  assign _zz_io_result_428 = ((_zz_io_result_426[0] && _zz_io_result_419[1]) ^ (_zz_io_result_419[0] && _zz_io_result_426[1]));
  always @(*) begin
    _zz_io_result_429[1] = ((_zz_io_result_426[0] && _zz_io_result_419[0]) ^ _zz_io_result_428);
    _zz_io_result_429[0] = ((_zz_io_result_426[1] && _zz_io_result_419[1]) ^ _zz_io_result_428);
  end

  assign _zz_io_result_430 = ((_zz_io_result_426[0] && _zz_io_result_420[1]) ^ (_zz_io_result_420[0] && _zz_io_result_426[1]));
  always @(*) begin
    _zz_io_result_431[1] = ((_zz_io_result_426[0] && _zz_io_result_420[0]) ^ _zz_io_result_430);
    _zz_io_result_431[0] = ((_zz_io_result_426[1] && _zz_io_result_420[1]) ^ _zz_io_result_430);
  end

  always @(*) begin
    _zz_io_result_418[3 : 2] = _zz_io_result_431;
    _zz_io_result_418[1 : 0] = _zz_io_result_429;
  end

  assign _zz_io_result_417 = _zz_io_result_418;
  assign _zz_io_result_433 = _zz_io_result_396[3 : 2];
  assign _zz_io_result_434 = _zz_io_result_396[1 : 0];
  assign _zz_io_result_435 = _zz_io_result_417[3 : 2];
  assign _zz_io_result_436 = _zz_io_result_417[1 : 0];
  assign _zz_io_result_437 = (_zz_io_result_433 ^ _zz_io_result_434);
  assign _zz_io_result_438 = (_zz_io_result_435 ^ _zz_io_result_436);
  assign _zz_io_result_440 = ((_zz_io_result_438[0] && _zz_io_result_437[1]) ^ (_zz_io_result_437[0] && _zz_io_result_438[1]));
  always @(*) begin
    _zz_io_result_441[1] = ((_zz_io_result_438[0] && _zz_io_result_437[0]) ^ _zz_io_result_440);
    _zz_io_result_441[0] = ((_zz_io_result_438[1] && _zz_io_result_437[1]) ^ _zz_io_result_440);
  end

  assign _zz_io_result_439 = _zz_io_result_441;
  always @(*) begin
    _zz_io_result_443[1] = _zz_io_result_439[0];
    _zz_io_result_443[0] = (_zz_io_result_439[0] ^ _zz_io_result_439[1]);
  end

  assign _zz_io_result_442 = _zz_io_result_443;
  assign _zz_io_result_444 = ((_zz_io_result_435[0] && _zz_io_result_433[1]) ^ (_zz_io_result_433[0] && _zz_io_result_435[1]));
  always @(*) begin
    _zz_io_result_445[1] = ((_zz_io_result_435[0] && _zz_io_result_433[0]) ^ _zz_io_result_444);
    _zz_io_result_445[0] = ((_zz_io_result_435[1] && _zz_io_result_433[1]) ^ _zz_io_result_444);
  end

  assign _zz_io_result_446 = ((_zz_io_result_436[0] && _zz_io_result_434[1]) ^ (_zz_io_result_434[0] && _zz_io_result_436[1]));
  always @(*) begin
    _zz_io_result_447[1] = ((_zz_io_result_436[0] && _zz_io_result_434[0]) ^ _zz_io_result_446);
    _zz_io_result_447[0] = ((_zz_io_result_436[1] && _zz_io_result_434[1]) ^ _zz_io_result_446);
  end

  always @(*) begin
    _zz_io_result_432[3 : 2] = (_zz_io_result_445 ^ _zz_io_result_442);
    _zz_io_result_432[1 : 0] = (_zz_io_result_447 ^ _zz_io_result_442);
  end

  assign _zz_io_result_449 = _zz_io_result_397[3 : 2];
  assign _zz_io_result_450 = _zz_io_result_397[1 : 0];
  assign _zz_io_result_451 = _zz_io_result_417[3 : 2];
  assign _zz_io_result_452 = _zz_io_result_417[1 : 0];
  assign _zz_io_result_453 = (_zz_io_result_449 ^ _zz_io_result_450);
  assign _zz_io_result_454 = (_zz_io_result_451 ^ _zz_io_result_452);
  assign _zz_io_result_456 = ((_zz_io_result_454[0] && _zz_io_result_453[1]) ^ (_zz_io_result_453[0] && _zz_io_result_454[1]));
  always @(*) begin
    _zz_io_result_457[1] = ((_zz_io_result_454[0] && _zz_io_result_453[0]) ^ _zz_io_result_456);
    _zz_io_result_457[0] = ((_zz_io_result_454[1] && _zz_io_result_453[1]) ^ _zz_io_result_456);
  end

  assign _zz_io_result_455 = _zz_io_result_457;
  always @(*) begin
    _zz_io_result_459[1] = _zz_io_result_455[0];
    _zz_io_result_459[0] = (_zz_io_result_455[0] ^ _zz_io_result_455[1]);
  end

  assign _zz_io_result_458 = _zz_io_result_459;
  assign _zz_io_result_460 = ((_zz_io_result_451[0] && _zz_io_result_449[1]) ^ (_zz_io_result_449[0] && _zz_io_result_451[1]));
  always @(*) begin
    _zz_io_result_461[1] = ((_zz_io_result_451[0] && _zz_io_result_449[0]) ^ _zz_io_result_460);
    _zz_io_result_461[0] = ((_zz_io_result_451[1] && _zz_io_result_449[1]) ^ _zz_io_result_460);
  end

  assign _zz_io_result_462 = ((_zz_io_result_452[0] && _zz_io_result_450[1]) ^ (_zz_io_result_450[0] && _zz_io_result_452[1]));
  always @(*) begin
    _zz_io_result_463[1] = ((_zz_io_result_452[0] && _zz_io_result_450[0]) ^ _zz_io_result_462);
    _zz_io_result_463[0] = ((_zz_io_result_452[1] && _zz_io_result_450[1]) ^ _zz_io_result_462);
  end

  always @(*) begin
    _zz_io_result_448[3 : 2] = (_zz_io_result_461 ^ _zz_io_result_458);
    _zz_io_result_448[1 : 0] = (_zz_io_result_463 ^ _zz_io_result_458);
  end

  always @(*) begin
    _zz_io_result_395[7 : 4] = _zz_io_result_448;
    _zz_io_result_395[3 : 0] = _zz_io_result_432;
  end

  assign _zz_io_result_394 = _zz_io_result_395;
  always @(*) begin
    _zz_io_result_465[7] = (_zz_io_result_394[5] ^ _zz_io_result_394[3]);
    _zz_io_result_465[6] = (_zz_io_result_394[7] ^ _zz_io_result_394[3]);
    _zz_io_result_465[5] = (_zz_io_result_394[6] ^ _zz_io_result_394[0]);
    _zz_io_result_465[4] = ((_zz_io_result_394[7] ^ _zz_io_result_394[5]) ^ _zz_io_result_394[3]);
    _zz_io_result_465[3] = ((((_zz_io_result_394[7] ^ _zz_io_result_394[6]) ^ _zz_io_result_394[5]) ^ _zz_io_result_394[4]) ^ _zz_io_result_394[3]);
    _zz_io_result_465[2] = ((((_zz_io_result_394[6] ^ _zz_io_result_394[5]) ^ _zz_io_result_394[3]) ^ _zz_io_result_394[2]) ^ _zz_io_result_394[0]);
    _zz_io_result_465[1] = ((_zz_io_result_394[5] ^ _zz_io_result_394[4]) ^ _zz_io_result_394[1]);
    _zz_io_result_465[0] = ((_zz_io_result_394[6] ^ _zz_io_result_394[4]) ^ _zz_io_result_394[1]);
  end

  assign _zz_io_result_464 = _zz_io_result_465;
  always @(*) begin
    _zz_io_result_391[7] = _zz_io_result_464[7];
    _zz_io_result_391[6] = (! _zz_io_result_464[6]);
    _zz_io_result_391[5] = (! _zz_io_result_464[5]);
    _zz_io_result_391[4] = _zz_io_result_464[4];
    _zz_io_result_391[3] = _zz_io_result_464[3];
    _zz_io_result_391[2] = _zz_io_result_464[2];
    _zz_io_result_391[1] = (! _zz_io_result_464[1]);
    _zz_io_result_391[0] = (! _zz_io_result_464[0]);
  end

  assign _zz_io_result_466 = _zz_io_result_1[23 : 16];
  always @(*) begin
    _zz_io_result_469[7] = (((((_zz_io_result_466[7] ^ _zz_io_result_466[6]) ^ _zz_io_result_466[5]) ^ _zz_io_result_466[2]) ^ _zz_io_result_466[1]) ^ _zz_io_result_466[0]);
    _zz_io_result_469[6] = (((_zz_io_result_466[6] ^ _zz_io_result_466[5]) ^ _zz_io_result_466[4]) ^ _zz_io_result_466[0]);
    _zz_io_result_469[5] = (((_zz_io_result_466[6] ^ _zz_io_result_466[5]) ^ _zz_io_result_466[1]) ^ _zz_io_result_466[0]);
    _zz_io_result_469[4] = (((_zz_io_result_466[7] ^ _zz_io_result_466[6]) ^ _zz_io_result_466[5]) ^ _zz_io_result_466[0]);
    _zz_io_result_469[3] = ((((_zz_io_result_466[7] ^ _zz_io_result_466[4]) ^ _zz_io_result_466[3]) ^ _zz_io_result_466[1]) ^ _zz_io_result_466[0]);
    _zz_io_result_469[2] = _zz_io_result_466[0];
    _zz_io_result_469[1] = ((_zz_io_result_466[6] ^ _zz_io_result_466[5]) ^ _zz_io_result_466[0]);
    _zz_io_result_469[0] = ((((_zz_io_result_466[6] ^ _zz_io_result_466[3]) ^ _zz_io_result_466[2]) ^ _zz_io_result_466[1]) ^ _zz_io_result_466[0]);
  end

  assign _zz_io_result_468 = _zz_io_result_469;
  assign _zz_io_result_472 = _zz_io_result_468[7 : 4];
  assign _zz_io_result_473 = _zz_io_result_468[3 : 0];
  assign _zz_io_result_474 = (_zz_io_result_472 ^ _zz_io_result_473);
  always @(*) begin
    _zz_io_result_475[3] = (_zz_io_result_474[2] ^ _zz_io_result_474[0]);
    _zz_io_result_475[2] = (_zz_io_result_474[3] ^ _zz_io_result_474[1]);
    _zz_io_result_475[1] = (_zz_io_result_474[1] ^ _zz_io_result_474[0]);
    _zz_io_result_475[0] = _zz_io_result_474[0];
  end

  assign _zz_io_result_477 = _zz_io_result_472[3 : 2];
  assign _zz_io_result_478 = _zz_io_result_472[1 : 0];
  assign _zz_io_result_479 = _zz_io_result_473[3 : 2];
  assign _zz_io_result_480 = _zz_io_result_473[1 : 0];
  assign _zz_io_result_481 = (_zz_io_result_477 ^ _zz_io_result_478);
  assign _zz_io_result_482 = (_zz_io_result_479 ^ _zz_io_result_480);
  assign _zz_io_result_484 = ((_zz_io_result_482[0] && _zz_io_result_481[1]) ^ (_zz_io_result_481[0] && _zz_io_result_482[1]));
  always @(*) begin
    _zz_io_result_485[1] = ((_zz_io_result_482[0] && _zz_io_result_481[0]) ^ _zz_io_result_484);
    _zz_io_result_485[0] = ((_zz_io_result_482[1] && _zz_io_result_481[1]) ^ _zz_io_result_484);
  end

  assign _zz_io_result_483 = _zz_io_result_485;
  always @(*) begin
    _zz_io_result_487[1] = _zz_io_result_483[0];
    _zz_io_result_487[0] = (_zz_io_result_483[0] ^ _zz_io_result_483[1]);
  end

  assign _zz_io_result_486 = _zz_io_result_487;
  assign _zz_io_result_488 = ((_zz_io_result_479[0] && _zz_io_result_477[1]) ^ (_zz_io_result_477[0] && _zz_io_result_479[1]));
  always @(*) begin
    _zz_io_result_489[1] = ((_zz_io_result_479[0] && _zz_io_result_477[0]) ^ _zz_io_result_488);
    _zz_io_result_489[0] = ((_zz_io_result_479[1] && _zz_io_result_477[1]) ^ _zz_io_result_488);
  end

  assign _zz_io_result_490 = ((_zz_io_result_480[0] && _zz_io_result_478[1]) ^ (_zz_io_result_478[0] && _zz_io_result_480[1]));
  always @(*) begin
    _zz_io_result_491[1] = ((_zz_io_result_480[0] && _zz_io_result_478[0]) ^ _zz_io_result_490);
    _zz_io_result_491[0] = ((_zz_io_result_480[1] && _zz_io_result_478[1]) ^ _zz_io_result_490);
  end

  always @(*) begin
    _zz_io_result_476[3 : 2] = (_zz_io_result_489 ^ _zz_io_result_486);
    _zz_io_result_476[1 : 0] = (_zz_io_result_491 ^ _zz_io_result_486);
  end

  assign _zz_io_result_492 = (_zz_io_result_475 ^ _zz_io_result_476);
  assign _zz_io_result_495 = _zz_io_result_492[3 : 2];
  assign _zz_io_result_496 = _zz_io_result_492[1 : 0];
  assign _zz_io_result_497 = (_zz_io_result_495 ^ _zz_io_result_496);
  always @(*) begin
    _zz_io_result_498[1] = _zz_io_result_497[1];
    _zz_io_result_498[0] = (_zz_io_result_497[0] ^ _zz_io_result_497[1]);
  end

  assign _zz_io_result_499 = ((_zz_io_result_496[0] && _zz_io_result_495[1]) ^ (_zz_io_result_495[0] && _zz_io_result_496[1]));
  always @(*) begin
    _zz_io_result_500[1] = ((_zz_io_result_496[0] && _zz_io_result_495[0]) ^ _zz_io_result_499);
    _zz_io_result_500[0] = ((_zz_io_result_496[1] && _zz_io_result_495[1]) ^ _zz_io_result_499);
  end

  assign _zz_io_result_501 = (_zz_io_result_498 ^ _zz_io_result_500);
  always @(*) begin
    _zz_io_result_503[1] = _zz_io_result_501[0];
    _zz_io_result_503[0] = _zz_io_result_501[1];
  end

  assign _zz_io_result_502 = _zz_io_result_503;
  assign _zz_io_result_504 = ((_zz_io_result_502[0] && _zz_io_result_495[1]) ^ (_zz_io_result_495[0] && _zz_io_result_502[1]));
  always @(*) begin
    _zz_io_result_505[1] = ((_zz_io_result_502[0] && _zz_io_result_495[0]) ^ _zz_io_result_504);
    _zz_io_result_505[0] = ((_zz_io_result_502[1] && _zz_io_result_495[1]) ^ _zz_io_result_504);
  end

  assign _zz_io_result_506 = ((_zz_io_result_502[0] && _zz_io_result_496[1]) ^ (_zz_io_result_496[0] && _zz_io_result_502[1]));
  always @(*) begin
    _zz_io_result_507[1] = ((_zz_io_result_502[0] && _zz_io_result_496[0]) ^ _zz_io_result_506);
    _zz_io_result_507[0] = ((_zz_io_result_502[1] && _zz_io_result_496[1]) ^ _zz_io_result_506);
  end

  always @(*) begin
    _zz_io_result_494[3 : 2] = _zz_io_result_507;
    _zz_io_result_494[1 : 0] = _zz_io_result_505;
  end

  assign _zz_io_result_493 = _zz_io_result_494;
  assign _zz_io_result_509 = _zz_io_result_472[3 : 2];
  assign _zz_io_result_510 = _zz_io_result_472[1 : 0];
  assign _zz_io_result_511 = _zz_io_result_493[3 : 2];
  assign _zz_io_result_512 = _zz_io_result_493[1 : 0];
  assign _zz_io_result_513 = (_zz_io_result_509 ^ _zz_io_result_510);
  assign _zz_io_result_514 = (_zz_io_result_511 ^ _zz_io_result_512);
  assign _zz_io_result_516 = ((_zz_io_result_514[0] && _zz_io_result_513[1]) ^ (_zz_io_result_513[0] && _zz_io_result_514[1]));
  always @(*) begin
    _zz_io_result_517[1] = ((_zz_io_result_514[0] && _zz_io_result_513[0]) ^ _zz_io_result_516);
    _zz_io_result_517[0] = ((_zz_io_result_514[1] && _zz_io_result_513[1]) ^ _zz_io_result_516);
  end

  assign _zz_io_result_515 = _zz_io_result_517;
  always @(*) begin
    _zz_io_result_519[1] = _zz_io_result_515[0];
    _zz_io_result_519[0] = (_zz_io_result_515[0] ^ _zz_io_result_515[1]);
  end

  assign _zz_io_result_518 = _zz_io_result_519;
  assign _zz_io_result_520 = ((_zz_io_result_511[0] && _zz_io_result_509[1]) ^ (_zz_io_result_509[0] && _zz_io_result_511[1]));
  always @(*) begin
    _zz_io_result_521[1] = ((_zz_io_result_511[0] && _zz_io_result_509[0]) ^ _zz_io_result_520);
    _zz_io_result_521[0] = ((_zz_io_result_511[1] && _zz_io_result_509[1]) ^ _zz_io_result_520);
  end

  assign _zz_io_result_522 = ((_zz_io_result_512[0] && _zz_io_result_510[1]) ^ (_zz_io_result_510[0] && _zz_io_result_512[1]));
  always @(*) begin
    _zz_io_result_523[1] = ((_zz_io_result_512[0] && _zz_io_result_510[0]) ^ _zz_io_result_522);
    _zz_io_result_523[0] = ((_zz_io_result_512[1] && _zz_io_result_510[1]) ^ _zz_io_result_522);
  end

  always @(*) begin
    _zz_io_result_508[3 : 2] = (_zz_io_result_521 ^ _zz_io_result_518);
    _zz_io_result_508[1 : 0] = (_zz_io_result_523 ^ _zz_io_result_518);
  end

  assign _zz_io_result_525 = _zz_io_result_473[3 : 2];
  assign _zz_io_result_526 = _zz_io_result_473[1 : 0];
  assign _zz_io_result_527 = _zz_io_result_493[3 : 2];
  assign _zz_io_result_528 = _zz_io_result_493[1 : 0];
  assign _zz_io_result_529 = (_zz_io_result_525 ^ _zz_io_result_526);
  assign _zz_io_result_530 = (_zz_io_result_527 ^ _zz_io_result_528);
  assign _zz_io_result_532 = ((_zz_io_result_530[0] && _zz_io_result_529[1]) ^ (_zz_io_result_529[0] && _zz_io_result_530[1]));
  always @(*) begin
    _zz_io_result_533[1] = ((_zz_io_result_530[0] && _zz_io_result_529[0]) ^ _zz_io_result_532);
    _zz_io_result_533[0] = ((_zz_io_result_530[1] && _zz_io_result_529[1]) ^ _zz_io_result_532);
  end

  assign _zz_io_result_531 = _zz_io_result_533;
  always @(*) begin
    _zz_io_result_535[1] = _zz_io_result_531[0];
    _zz_io_result_535[0] = (_zz_io_result_531[0] ^ _zz_io_result_531[1]);
  end

  assign _zz_io_result_534 = _zz_io_result_535;
  assign _zz_io_result_536 = ((_zz_io_result_527[0] && _zz_io_result_525[1]) ^ (_zz_io_result_525[0] && _zz_io_result_527[1]));
  always @(*) begin
    _zz_io_result_537[1] = ((_zz_io_result_527[0] && _zz_io_result_525[0]) ^ _zz_io_result_536);
    _zz_io_result_537[0] = ((_zz_io_result_527[1] && _zz_io_result_525[1]) ^ _zz_io_result_536);
  end

  assign _zz_io_result_538 = ((_zz_io_result_528[0] && _zz_io_result_526[1]) ^ (_zz_io_result_526[0] && _zz_io_result_528[1]));
  always @(*) begin
    _zz_io_result_539[1] = ((_zz_io_result_528[0] && _zz_io_result_526[0]) ^ _zz_io_result_538);
    _zz_io_result_539[0] = ((_zz_io_result_528[1] && _zz_io_result_526[1]) ^ _zz_io_result_538);
  end

  always @(*) begin
    _zz_io_result_524[3 : 2] = (_zz_io_result_537 ^ _zz_io_result_534);
    _zz_io_result_524[1 : 0] = (_zz_io_result_539 ^ _zz_io_result_534);
  end

  always @(*) begin
    _zz_io_result_471[7 : 4] = _zz_io_result_524;
    _zz_io_result_471[3 : 0] = _zz_io_result_508;
  end

  assign _zz_io_result_470 = _zz_io_result_471;
  always @(*) begin
    _zz_io_result_541[7] = (_zz_io_result_470[5] ^ _zz_io_result_470[3]);
    _zz_io_result_541[6] = (_zz_io_result_470[7] ^ _zz_io_result_470[3]);
    _zz_io_result_541[5] = (_zz_io_result_470[6] ^ _zz_io_result_470[0]);
    _zz_io_result_541[4] = ((_zz_io_result_470[7] ^ _zz_io_result_470[5]) ^ _zz_io_result_470[3]);
    _zz_io_result_541[3] = ((((_zz_io_result_470[7] ^ _zz_io_result_470[6]) ^ _zz_io_result_470[5]) ^ _zz_io_result_470[4]) ^ _zz_io_result_470[3]);
    _zz_io_result_541[2] = ((((_zz_io_result_470[6] ^ _zz_io_result_470[5]) ^ _zz_io_result_470[3]) ^ _zz_io_result_470[2]) ^ _zz_io_result_470[0]);
    _zz_io_result_541[1] = ((_zz_io_result_470[5] ^ _zz_io_result_470[4]) ^ _zz_io_result_470[1]);
    _zz_io_result_541[0] = ((_zz_io_result_470[6] ^ _zz_io_result_470[4]) ^ _zz_io_result_470[1]);
  end

  assign _zz_io_result_540 = _zz_io_result_541;
  always @(*) begin
    _zz_io_result_467[7] = _zz_io_result_540[7];
    _zz_io_result_467[6] = (! _zz_io_result_540[6]);
    _zz_io_result_467[5] = (! _zz_io_result_540[5]);
    _zz_io_result_467[4] = _zz_io_result_540[4];
    _zz_io_result_467[3] = _zz_io_result_540[3];
    _zz_io_result_467[2] = _zz_io_result_540[2];
    _zz_io_result_467[1] = (! _zz_io_result_540[1]);
    _zz_io_result_467[0] = (! _zz_io_result_540[0]);
  end

  assign _zz_io_result_542 = _zz_io_result_1[31 : 24];
  always @(*) begin
    _zz_io_result_545[7] = (((((_zz_io_result_542[7] ^ _zz_io_result_542[6]) ^ _zz_io_result_542[5]) ^ _zz_io_result_542[2]) ^ _zz_io_result_542[1]) ^ _zz_io_result_542[0]);
    _zz_io_result_545[6] = (((_zz_io_result_542[6] ^ _zz_io_result_542[5]) ^ _zz_io_result_542[4]) ^ _zz_io_result_542[0]);
    _zz_io_result_545[5] = (((_zz_io_result_542[6] ^ _zz_io_result_542[5]) ^ _zz_io_result_542[1]) ^ _zz_io_result_542[0]);
    _zz_io_result_545[4] = (((_zz_io_result_542[7] ^ _zz_io_result_542[6]) ^ _zz_io_result_542[5]) ^ _zz_io_result_542[0]);
    _zz_io_result_545[3] = ((((_zz_io_result_542[7] ^ _zz_io_result_542[4]) ^ _zz_io_result_542[3]) ^ _zz_io_result_542[1]) ^ _zz_io_result_542[0]);
    _zz_io_result_545[2] = _zz_io_result_542[0];
    _zz_io_result_545[1] = ((_zz_io_result_542[6] ^ _zz_io_result_542[5]) ^ _zz_io_result_542[0]);
    _zz_io_result_545[0] = ((((_zz_io_result_542[6] ^ _zz_io_result_542[3]) ^ _zz_io_result_542[2]) ^ _zz_io_result_542[1]) ^ _zz_io_result_542[0]);
  end

  assign _zz_io_result_544 = _zz_io_result_545;
  assign _zz_io_result_548 = _zz_io_result_544[7 : 4];
  assign _zz_io_result_549 = _zz_io_result_544[3 : 0];
  assign _zz_io_result_550 = (_zz_io_result_548 ^ _zz_io_result_549);
  always @(*) begin
    _zz_io_result_551[3] = (_zz_io_result_550[2] ^ _zz_io_result_550[0]);
    _zz_io_result_551[2] = (_zz_io_result_550[3] ^ _zz_io_result_550[1]);
    _zz_io_result_551[1] = (_zz_io_result_550[1] ^ _zz_io_result_550[0]);
    _zz_io_result_551[0] = _zz_io_result_550[0];
  end

  assign _zz_io_result_553 = _zz_io_result_548[3 : 2];
  assign _zz_io_result_554 = _zz_io_result_548[1 : 0];
  assign _zz_io_result_555 = _zz_io_result_549[3 : 2];
  assign _zz_io_result_556 = _zz_io_result_549[1 : 0];
  assign _zz_io_result_557 = (_zz_io_result_553 ^ _zz_io_result_554);
  assign _zz_io_result_558 = (_zz_io_result_555 ^ _zz_io_result_556);
  assign _zz_io_result_560 = ((_zz_io_result_558[0] && _zz_io_result_557[1]) ^ (_zz_io_result_557[0] && _zz_io_result_558[1]));
  always @(*) begin
    _zz_io_result_561[1] = ((_zz_io_result_558[0] && _zz_io_result_557[0]) ^ _zz_io_result_560);
    _zz_io_result_561[0] = ((_zz_io_result_558[1] && _zz_io_result_557[1]) ^ _zz_io_result_560);
  end

  assign _zz_io_result_559 = _zz_io_result_561;
  always @(*) begin
    _zz_io_result_563[1] = _zz_io_result_559[0];
    _zz_io_result_563[0] = (_zz_io_result_559[0] ^ _zz_io_result_559[1]);
  end

  assign _zz_io_result_562 = _zz_io_result_563;
  assign _zz_io_result_564 = ((_zz_io_result_555[0] && _zz_io_result_553[1]) ^ (_zz_io_result_553[0] && _zz_io_result_555[1]));
  always @(*) begin
    _zz_io_result_565[1] = ((_zz_io_result_555[0] && _zz_io_result_553[0]) ^ _zz_io_result_564);
    _zz_io_result_565[0] = ((_zz_io_result_555[1] && _zz_io_result_553[1]) ^ _zz_io_result_564);
  end

  assign _zz_io_result_566 = ((_zz_io_result_556[0] && _zz_io_result_554[1]) ^ (_zz_io_result_554[0] && _zz_io_result_556[1]));
  always @(*) begin
    _zz_io_result_567[1] = ((_zz_io_result_556[0] && _zz_io_result_554[0]) ^ _zz_io_result_566);
    _zz_io_result_567[0] = ((_zz_io_result_556[1] && _zz_io_result_554[1]) ^ _zz_io_result_566);
  end

  always @(*) begin
    _zz_io_result_552[3 : 2] = (_zz_io_result_565 ^ _zz_io_result_562);
    _zz_io_result_552[1 : 0] = (_zz_io_result_567 ^ _zz_io_result_562);
  end

  assign _zz_io_result_568 = (_zz_io_result_551 ^ _zz_io_result_552);
  assign _zz_io_result_571 = _zz_io_result_568[3 : 2];
  assign _zz_io_result_572 = _zz_io_result_568[1 : 0];
  assign _zz_io_result_573 = (_zz_io_result_571 ^ _zz_io_result_572);
  always @(*) begin
    _zz_io_result_574[1] = _zz_io_result_573[1];
    _zz_io_result_574[0] = (_zz_io_result_573[0] ^ _zz_io_result_573[1]);
  end

  assign _zz_io_result_575 = ((_zz_io_result_572[0] && _zz_io_result_571[1]) ^ (_zz_io_result_571[0] && _zz_io_result_572[1]));
  always @(*) begin
    _zz_io_result_576[1] = ((_zz_io_result_572[0] && _zz_io_result_571[0]) ^ _zz_io_result_575);
    _zz_io_result_576[0] = ((_zz_io_result_572[1] && _zz_io_result_571[1]) ^ _zz_io_result_575);
  end

  assign _zz_io_result_577 = (_zz_io_result_574 ^ _zz_io_result_576);
  always @(*) begin
    _zz_io_result_579[1] = _zz_io_result_577[0];
    _zz_io_result_579[0] = _zz_io_result_577[1];
  end

  assign _zz_io_result_578 = _zz_io_result_579;
  assign _zz_io_result_580 = ((_zz_io_result_578[0] && _zz_io_result_571[1]) ^ (_zz_io_result_571[0] && _zz_io_result_578[1]));
  always @(*) begin
    _zz_io_result_581[1] = ((_zz_io_result_578[0] && _zz_io_result_571[0]) ^ _zz_io_result_580);
    _zz_io_result_581[0] = ((_zz_io_result_578[1] && _zz_io_result_571[1]) ^ _zz_io_result_580);
  end

  assign _zz_io_result_582 = ((_zz_io_result_578[0] && _zz_io_result_572[1]) ^ (_zz_io_result_572[0] && _zz_io_result_578[1]));
  always @(*) begin
    _zz_io_result_583[1] = ((_zz_io_result_578[0] && _zz_io_result_572[0]) ^ _zz_io_result_582);
    _zz_io_result_583[0] = ((_zz_io_result_578[1] && _zz_io_result_572[1]) ^ _zz_io_result_582);
  end

  always @(*) begin
    _zz_io_result_570[3 : 2] = _zz_io_result_583;
    _zz_io_result_570[1 : 0] = _zz_io_result_581;
  end

  assign _zz_io_result_569 = _zz_io_result_570;
  assign _zz_io_result_585 = _zz_io_result_548[3 : 2];
  assign _zz_io_result_586 = _zz_io_result_548[1 : 0];
  assign _zz_io_result_587 = _zz_io_result_569[3 : 2];
  assign _zz_io_result_588 = _zz_io_result_569[1 : 0];
  assign _zz_io_result_589 = (_zz_io_result_585 ^ _zz_io_result_586);
  assign _zz_io_result_590 = (_zz_io_result_587 ^ _zz_io_result_588);
  assign _zz_io_result_592 = ((_zz_io_result_590[0] && _zz_io_result_589[1]) ^ (_zz_io_result_589[0] && _zz_io_result_590[1]));
  always @(*) begin
    _zz_io_result_593[1] = ((_zz_io_result_590[0] && _zz_io_result_589[0]) ^ _zz_io_result_592);
    _zz_io_result_593[0] = ((_zz_io_result_590[1] && _zz_io_result_589[1]) ^ _zz_io_result_592);
  end

  assign _zz_io_result_591 = _zz_io_result_593;
  always @(*) begin
    _zz_io_result_595[1] = _zz_io_result_591[0];
    _zz_io_result_595[0] = (_zz_io_result_591[0] ^ _zz_io_result_591[1]);
  end

  assign _zz_io_result_594 = _zz_io_result_595;
  assign _zz_io_result_596 = ((_zz_io_result_587[0] && _zz_io_result_585[1]) ^ (_zz_io_result_585[0] && _zz_io_result_587[1]));
  always @(*) begin
    _zz_io_result_597[1] = ((_zz_io_result_587[0] && _zz_io_result_585[0]) ^ _zz_io_result_596);
    _zz_io_result_597[0] = ((_zz_io_result_587[1] && _zz_io_result_585[1]) ^ _zz_io_result_596);
  end

  assign _zz_io_result_598 = ((_zz_io_result_588[0] && _zz_io_result_586[1]) ^ (_zz_io_result_586[0] && _zz_io_result_588[1]));
  always @(*) begin
    _zz_io_result_599[1] = ((_zz_io_result_588[0] && _zz_io_result_586[0]) ^ _zz_io_result_598);
    _zz_io_result_599[0] = ((_zz_io_result_588[1] && _zz_io_result_586[1]) ^ _zz_io_result_598);
  end

  always @(*) begin
    _zz_io_result_584[3 : 2] = (_zz_io_result_597 ^ _zz_io_result_594);
    _zz_io_result_584[1 : 0] = (_zz_io_result_599 ^ _zz_io_result_594);
  end

  assign _zz_io_result_601 = _zz_io_result_549[3 : 2];
  assign _zz_io_result_602 = _zz_io_result_549[1 : 0];
  assign _zz_io_result_603 = _zz_io_result_569[3 : 2];
  assign _zz_io_result_604 = _zz_io_result_569[1 : 0];
  assign _zz_io_result_605 = (_zz_io_result_601 ^ _zz_io_result_602);
  assign _zz_io_result_606 = (_zz_io_result_603 ^ _zz_io_result_604);
  assign _zz_io_result_608 = ((_zz_io_result_606[0] && _zz_io_result_605[1]) ^ (_zz_io_result_605[0] && _zz_io_result_606[1]));
  always @(*) begin
    _zz_io_result_609[1] = ((_zz_io_result_606[0] && _zz_io_result_605[0]) ^ _zz_io_result_608);
    _zz_io_result_609[0] = ((_zz_io_result_606[1] && _zz_io_result_605[1]) ^ _zz_io_result_608);
  end

  assign _zz_io_result_607 = _zz_io_result_609;
  always @(*) begin
    _zz_io_result_611[1] = _zz_io_result_607[0];
    _zz_io_result_611[0] = (_zz_io_result_607[0] ^ _zz_io_result_607[1]);
  end

  assign _zz_io_result_610 = _zz_io_result_611;
  assign _zz_io_result_612 = ((_zz_io_result_603[0] && _zz_io_result_601[1]) ^ (_zz_io_result_601[0] && _zz_io_result_603[1]));
  always @(*) begin
    _zz_io_result_613[1] = ((_zz_io_result_603[0] && _zz_io_result_601[0]) ^ _zz_io_result_612);
    _zz_io_result_613[0] = ((_zz_io_result_603[1] && _zz_io_result_601[1]) ^ _zz_io_result_612);
  end

  assign _zz_io_result_614 = ((_zz_io_result_604[0] && _zz_io_result_602[1]) ^ (_zz_io_result_602[0] && _zz_io_result_604[1]));
  always @(*) begin
    _zz_io_result_615[1] = ((_zz_io_result_604[0] && _zz_io_result_602[0]) ^ _zz_io_result_614);
    _zz_io_result_615[0] = ((_zz_io_result_604[1] && _zz_io_result_602[1]) ^ _zz_io_result_614);
  end

  always @(*) begin
    _zz_io_result_600[3 : 2] = (_zz_io_result_613 ^ _zz_io_result_610);
    _zz_io_result_600[1 : 0] = (_zz_io_result_615 ^ _zz_io_result_610);
  end

  always @(*) begin
    _zz_io_result_547[7 : 4] = _zz_io_result_600;
    _zz_io_result_547[3 : 0] = _zz_io_result_584;
  end

  assign _zz_io_result_546 = _zz_io_result_547;
  always @(*) begin
    _zz_io_result_617[7] = (_zz_io_result_546[5] ^ _zz_io_result_546[3]);
    _zz_io_result_617[6] = (_zz_io_result_546[7] ^ _zz_io_result_546[3]);
    _zz_io_result_617[5] = (_zz_io_result_546[6] ^ _zz_io_result_546[0]);
    _zz_io_result_617[4] = ((_zz_io_result_546[7] ^ _zz_io_result_546[5]) ^ _zz_io_result_546[3]);
    _zz_io_result_617[3] = ((((_zz_io_result_546[7] ^ _zz_io_result_546[6]) ^ _zz_io_result_546[5]) ^ _zz_io_result_546[4]) ^ _zz_io_result_546[3]);
    _zz_io_result_617[2] = ((((_zz_io_result_546[6] ^ _zz_io_result_546[5]) ^ _zz_io_result_546[3]) ^ _zz_io_result_546[2]) ^ _zz_io_result_546[0]);
    _zz_io_result_617[1] = ((_zz_io_result_546[5] ^ _zz_io_result_546[4]) ^ _zz_io_result_546[1]);
    _zz_io_result_617[0] = ((_zz_io_result_546[6] ^ _zz_io_result_546[4]) ^ _zz_io_result_546[1]);
  end

  assign _zz_io_result_616 = _zz_io_result_617;
  always @(*) begin
    _zz_io_result_543[7] = _zz_io_result_616[7];
    _zz_io_result_543[6] = (! _zz_io_result_616[6]);
    _zz_io_result_543[5] = (! _zz_io_result_616[5]);
    _zz_io_result_543[4] = _zz_io_result_616[4];
    _zz_io_result_543[3] = _zz_io_result_616[3];
    _zz_io_result_543[2] = _zz_io_result_616[2];
    _zz_io_result_543[1] = (! _zz_io_result_616[1]);
    _zz_io_result_543[0] = (! _zz_io_result_616[0]);
  end

  assign _zz_io_result_619 = _zz_io_result_2[7 : 0];
  always @(*) begin
    _zz_io_result_622[7] = (((((_zz_io_result_619[7] ^ _zz_io_result_619[6]) ^ _zz_io_result_619[5]) ^ _zz_io_result_619[2]) ^ _zz_io_result_619[1]) ^ _zz_io_result_619[0]);
    _zz_io_result_622[6] = (((_zz_io_result_619[6] ^ _zz_io_result_619[5]) ^ _zz_io_result_619[4]) ^ _zz_io_result_619[0]);
    _zz_io_result_622[5] = (((_zz_io_result_619[6] ^ _zz_io_result_619[5]) ^ _zz_io_result_619[1]) ^ _zz_io_result_619[0]);
    _zz_io_result_622[4] = (((_zz_io_result_619[7] ^ _zz_io_result_619[6]) ^ _zz_io_result_619[5]) ^ _zz_io_result_619[0]);
    _zz_io_result_622[3] = ((((_zz_io_result_619[7] ^ _zz_io_result_619[4]) ^ _zz_io_result_619[3]) ^ _zz_io_result_619[1]) ^ _zz_io_result_619[0]);
    _zz_io_result_622[2] = _zz_io_result_619[0];
    _zz_io_result_622[1] = ((_zz_io_result_619[6] ^ _zz_io_result_619[5]) ^ _zz_io_result_619[0]);
    _zz_io_result_622[0] = ((((_zz_io_result_619[6] ^ _zz_io_result_619[3]) ^ _zz_io_result_619[2]) ^ _zz_io_result_619[1]) ^ _zz_io_result_619[0]);
  end

  assign _zz_io_result_621 = _zz_io_result_622;
  assign _zz_io_result_625 = _zz_io_result_621[7 : 4];
  assign _zz_io_result_626 = _zz_io_result_621[3 : 0];
  assign _zz_io_result_627 = (_zz_io_result_625 ^ _zz_io_result_626);
  always @(*) begin
    _zz_io_result_628[3] = (_zz_io_result_627[2] ^ _zz_io_result_627[0]);
    _zz_io_result_628[2] = (_zz_io_result_627[3] ^ _zz_io_result_627[1]);
    _zz_io_result_628[1] = (_zz_io_result_627[1] ^ _zz_io_result_627[0]);
    _zz_io_result_628[0] = _zz_io_result_627[0];
  end

  assign _zz_io_result_630 = _zz_io_result_625[3 : 2];
  assign _zz_io_result_631 = _zz_io_result_625[1 : 0];
  assign _zz_io_result_632 = _zz_io_result_626[3 : 2];
  assign _zz_io_result_633 = _zz_io_result_626[1 : 0];
  assign _zz_io_result_634 = (_zz_io_result_630 ^ _zz_io_result_631);
  assign _zz_io_result_635 = (_zz_io_result_632 ^ _zz_io_result_633);
  assign _zz_io_result_637 = ((_zz_io_result_635[0] && _zz_io_result_634[1]) ^ (_zz_io_result_634[0] && _zz_io_result_635[1]));
  always @(*) begin
    _zz_io_result_638[1] = ((_zz_io_result_635[0] && _zz_io_result_634[0]) ^ _zz_io_result_637);
    _zz_io_result_638[0] = ((_zz_io_result_635[1] && _zz_io_result_634[1]) ^ _zz_io_result_637);
  end

  assign _zz_io_result_636 = _zz_io_result_638;
  always @(*) begin
    _zz_io_result_640[1] = _zz_io_result_636[0];
    _zz_io_result_640[0] = (_zz_io_result_636[0] ^ _zz_io_result_636[1]);
  end

  assign _zz_io_result_639 = _zz_io_result_640;
  assign _zz_io_result_641 = ((_zz_io_result_632[0] && _zz_io_result_630[1]) ^ (_zz_io_result_630[0] && _zz_io_result_632[1]));
  always @(*) begin
    _zz_io_result_642[1] = ((_zz_io_result_632[0] && _zz_io_result_630[0]) ^ _zz_io_result_641);
    _zz_io_result_642[0] = ((_zz_io_result_632[1] && _zz_io_result_630[1]) ^ _zz_io_result_641);
  end

  assign _zz_io_result_643 = ((_zz_io_result_633[0] && _zz_io_result_631[1]) ^ (_zz_io_result_631[0] && _zz_io_result_633[1]));
  always @(*) begin
    _zz_io_result_644[1] = ((_zz_io_result_633[0] && _zz_io_result_631[0]) ^ _zz_io_result_643);
    _zz_io_result_644[0] = ((_zz_io_result_633[1] && _zz_io_result_631[1]) ^ _zz_io_result_643);
  end

  always @(*) begin
    _zz_io_result_629[3 : 2] = (_zz_io_result_642 ^ _zz_io_result_639);
    _zz_io_result_629[1 : 0] = (_zz_io_result_644 ^ _zz_io_result_639);
  end

  assign _zz_io_result_645 = (_zz_io_result_628 ^ _zz_io_result_629);
  assign _zz_io_result_648 = _zz_io_result_645[3 : 2];
  assign _zz_io_result_649 = _zz_io_result_645[1 : 0];
  assign _zz_io_result_650 = (_zz_io_result_648 ^ _zz_io_result_649);
  always @(*) begin
    _zz_io_result_651[1] = _zz_io_result_650[1];
    _zz_io_result_651[0] = (_zz_io_result_650[0] ^ _zz_io_result_650[1]);
  end

  assign _zz_io_result_652 = ((_zz_io_result_649[0] && _zz_io_result_648[1]) ^ (_zz_io_result_648[0] && _zz_io_result_649[1]));
  always @(*) begin
    _zz_io_result_653[1] = ((_zz_io_result_649[0] && _zz_io_result_648[0]) ^ _zz_io_result_652);
    _zz_io_result_653[0] = ((_zz_io_result_649[1] && _zz_io_result_648[1]) ^ _zz_io_result_652);
  end

  assign _zz_io_result_654 = (_zz_io_result_651 ^ _zz_io_result_653);
  always @(*) begin
    _zz_io_result_656[1] = _zz_io_result_654[0];
    _zz_io_result_656[0] = _zz_io_result_654[1];
  end

  assign _zz_io_result_655 = _zz_io_result_656;
  assign _zz_io_result_657 = ((_zz_io_result_655[0] && _zz_io_result_648[1]) ^ (_zz_io_result_648[0] && _zz_io_result_655[1]));
  always @(*) begin
    _zz_io_result_658[1] = ((_zz_io_result_655[0] && _zz_io_result_648[0]) ^ _zz_io_result_657);
    _zz_io_result_658[0] = ((_zz_io_result_655[1] && _zz_io_result_648[1]) ^ _zz_io_result_657);
  end

  assign _zz_io_result_659 = ((_zz_io_result_655[0] && _zz_io_result_649[1]) ^ (_zz_io_result_649[0] && _zz_io_result_655[1]));
  always @(*) begin
    _zz_io_result_660[1] = ((_zz_io_result_655[0] && _zz_io_result_649[0]) ^ _zz_io_result_659);
    _zz_io_result_660[0] = ((_zz_io_result_655[1] && _zz_io_result_649[1]) ^ _zz_io_result_659);
  end

  always @(*) begin
    _zz_io_result_647[3 : 2] = _zz_io_result_660;
    _zz_io_result_647[1 : 0] = _zz_io_result_658;
  end

  assign _zz_io_result_646 = _zz_io_result_647;
  assign _zz_io_result_662 = _zz_io_result_625[3 : 2];
  assign _zz_io_result_663 = _zz_io_result_625[1 : 0];
  assign _zz_io_result_664 = _zz_io_result_646[3 : 2];
  assign _zz_io_result_665 = _zz_io_result_646[1 : 0];
  assign _zz_io_result_666 = (_zz_io_result_662 ^ _zz_io_result_663);
  assign _zz_io_result_667 = (_zz_io_result_664 ^ _zz_io_result_665);
  assign _zz_io_result_669 = ((_zz_io_result_667[0] && _zz_io_result_666[1]) ^ (_zz_io_result_666[0] && _zz_io_result_667[1]));
  always @(*) begin
    _zz_io_result_670[1] = ((_zz_io_result_667[0] && _zz_io_result_666[0]) ^ _zz_io_result_669);
    _zz_io_result_670[0] = ((_zz_io_result_667[1] && _zz_io_result_666[1]) ^ _zz_io_result_669);
  end

  assign _zz_io_result_668 = _zz_io_result_670;
  always @(*) begin
    _zz_io_result_672[1] = _zz_io_result_668[0];
    _zz_io_result_672[0] = (_zz_io_result_668[0] ^ _zz_io_result_668[1]);
  end

  assign _zz_io_result_671 = _zz_io_result_672;
  assign _zz_io_result_673 = ((_zz_io_result_664[0] && _zz_io_result_662[1]) ^ (_zz_io_result_662[0] && _zz_io_result_664[1]));
  always @(*) begin
    _zz_io_result_674[1] = ((_zz_io_result_664[0] && _zz_io_result_662[0]) ^ _zz_io_result_673);
    _zz_io_result_674[0] = ((_zz_io_result_664[1] && _zz_io_result_662[1]) ^ _zz_io_result_673);
  end

  assign _zz_io_result_675 = ((_zz_io_result_665[0] && _zz_io_result_663[1]) ^ (_zz_io_result_663[0] && _zz_io_result_665[1]));
  always @(*) begin
    _zz_io_result_676[1] = ((_zz_io_result_665[0] && _zz_io_result_663[0]) ^ _zz_io_result_675);
    _zz_io_result_676[0] = ((_zz_io_result_665[1] && _zz_io_result_663[1]) ^ _zz_io_result_675);
  end

  always @(*) begin
    _zz_io_result_661[3 : 2] = (_zz_io_result_674 ^ _zz_io_result_671);
    _zz_io_result_661[1 : 0] = (_zz_io_result_676 ^ _zz_io_result_671);
  end

  assign _zz_io_result_678 = _zz_io_result_626[3 : 2];
  assign _zz_io_result_679 = _zz_io_result_626[1 : 0];
  assign _zz_io_result_680 = _zz_io_result_646[3 : 2];
  assign _zz_io_result_681 = _zz_io_result_646[1 : 0];
  assign _zz_io_result_682 = (_zz_io_result_678 ^ _zz_io_result_679);
  assign _zz_io_result_683 = (_zz_io_result_680 ^ _zz_io_result_681);
  assign _zz_io_result_685 = ((_zz_io_result_683[0] && _zz_io_result_682[1]) ^ (_zz_io_result_682[0] && _zz_io_result_683[1]));
  always @(*) begin
    _zz_io_result_686[1] = ((_zz_io_result_683[0] && _zz_io_result_682[0]) ^ _zz_io_result_685);
    _zz_io_result_686[0] = ((_zz_io_result_683[1] && _zz_io_result_682[1]) ^ _zz_io_result_685);
  end

  assign _zz_io_result_684 = _zz_io_result_686;
  always @(*) begin
    _zz_io_result_688[1] = _zz_io_result_684[0];
    _zz_io_result_688[0] = (_zz_io_result_684[0] ^ _zz_io_result_684[1]);
  end

  assign _zz_io_result_687 = _zz_io_result_688;
  assign _zz_io_result_689 = ((_zz_io_result_680[0] && _zz_io_result_678[1]) ^ (_zz_io_result_678[0] && _zz_io_result_680[1]));
  always @(*) begin
    _zz_io_result_690[1] = ((_zz_io_result_680[0] && _zz_io_result_678[0]) ^ _zz_io_result_689);
    _zz_io_result_690[0] = ((_zz_io_result_680[1] && _zz_io_result_678[1]) ^ _zz_io_result_689);
  end

  assign _zz_io_result_691 = ((_zz_io_result_681[0] && _zz_io_result_679[1]) ^ (_zz_io_result_679[0] && _zz_io_result_681[1]));
  always @(*) begin
    _zz_io_result_692[1] = ((_zz_io_result_681[0] && _zz_io_result_679[0]) ^ _zz_io_result_691);
    _zz_io_result_692[0] = ((_zz_io_result_681[1] && _zz_io_result_679[1]) ^ _zz_io_result_691);
  end

  always @(*) begin
    _zz_io_result_677[3 : 2] = (_zz_io_result_690 ^ _zz_io_result_687);
    _zz_io_result_677[1 : 0] = (_zz_io_result_692 ^ _zz_io_result_687);
  end

  always @(*) begin
    _zz_io_result_624[7 : 4] = _zz_io_result_677;
    _zz_io_result_624[3 : 0] = _zz_io_result_661;
  end

  assign _zz_io_result_623 = _zz_io_result_624;
  always @(*) begin
    _zz_io_result_694[7] = (_zz_io_result_623[5] ^ _zz_io_result_623[3]);
    _zz_io_result_694[6] = (_zz_io_result_623[7] ^ _zz_io_result_623[3]);
    _zz_io_result_694[5] = (_zz_io_result_623[6] ^ _zz_io_result_623[0]);
    _zz_io_result_694[4] = ((_zz_io_result_623[7] ^ _zz_io_result_623[5]) ^ _zz_io_result_623[3]);
    _zz_io_result_694[3] = ((((_zz_io_result_623[7] ^ _zz_io_result_623[6]) ^ _zz_io_result_623[5]) ^ _zz_io_result_623[4]) ^ _zz_io_result_623[3]);
    _zz_io_result_694[2] = ((((_zz_io_result_623[6] ^ _zz_io_result_623[5]) ^ _zz_io_result_623[3]) ^ _zz_io_result_623[2]) ^ _zz_io_result_623[0]);
    _zz_io_result_694[1] = ((_zz_io_result_623[5] ^ _zz_io_result_623[4]) ^ _zz_io_result_623[1]);
    _zz_io_result_694[0] = ((_zz_io_result_623[6] ^ _zz_io_result_623[4]) ^ _zz_io_result_623[1]);
  end

  assign _zz_io_result_693 = _zz_io_result_694;
  always @(*) begin
    _zz_io_result_620[7] = _zz_io_result_693[7];
    _zz_io_result_620[6] = (! _zz_io_result_693[6]);
    _zz_io_result_620[5] = (! _zz_io_result_693[5]);
    _zz_io_result_620[4] = _zz_io_result_693[4];
    _zz_io_result_620[3] = _zz_io_result_693[3];
    _zz_io_result_620[2] = _zz_io_result_693[2];
    _zz_io_result_620[1] = (! _zz_io_result_693[1]);
    _zz_io_result_620[0] = (! _zz_io_result_693[0]);
  end

  always @(*) begin
    _zz_io_result_618[7 : 0] = _zz_io_result_620;
    _zz_io_result_618[15 : 8] = _zz_io_result_696;
    _zz_io_result_618[23 : 16] = _zz_io_result_772;
    _zz_io_result_618[31 : 24] = _zz_io_result_848;
  end

  assign _zz_io_result_695 = _zz_io_result_2[15 : 8];
  always @(*) begin
    _zz_io_result_698[7] = (((((_zz_io_result_695[7] ^ _zz_io_result_695[6]) ^ _zz_io_result_695[5]) ^ _zz_io_result_695[2]) ^ _zz_io_result_695[1]) ^ _zz_io_result_695[0]);
    _zz_io_result_698[6] = (((_zz_io_result_695[6] ^ _zz_io_result_695[5]) ^ _zz_io_result_695[4]) ^ _zz_io_result_695[0]);
    _zz_io_result_698[5] = (((_zz_io_result_695[6] ^ _zz_io_result_695[5]) ^ _zz_io_result_695[1]) ^ _zz_io_result_695[0]);
    _zz_io_result_698[4] = (((_zz_io_result_695[7] ^ _zz_io_result_695[6]) ^ _zz_io_result_695[5]) ^ _zz_io_result_695[0]);
    _zz_io_result_698[3] = ((((_zz_io_result_695[7] ^ _zz_io_result_695[4]) ^ _zz_io_result_695[3]) ^ _zz_io_result_695[1]) ^ _zz_io_result_695[0]);
    _zz_io_result_698[2] = _zz_io_result_695[0];
    _zz_io_result_698[1] = ((_zz_io_result_695[6] ^ _zz_io_result_695[5]) ^ _zz_io_result_695[0]);
    _zz_io_result_698[0] = ((((_zz_io_result_695[6] ^ _zz_io_result_695[3]) ^ _zz_io_result_695[2]) ^ _zz_io_result_695[1]) ^ _zz_io_result_695[0]);
  end

  assign _zz_io_result_697 = _zz_io_result_698;
  assign _zz_io_result_701 = _zz_io_result_697[7 : 4];
  assign _zz_io_result_702 = _zz_io_result_697[3 : 0];
  assign _zz_io_result_703 = (_zz_io_result_701 ^ _zz_io_result_702);
  always @(*) begin
    _zz_io_result_704[3] = (_zz_io_result_703[2] ^ _zz_io_result_703[0]);
    _zz_io_result_704[2] = (_zz_io_result_703[3] ^ _zz_io_result_703[1]);
    _zz_io_result_704[1] = (_zz_io_result_703[1] ^ _zz_io_result_703[0]);
    _zz_io_result_704[0] = _zz_io_result_703[0];
  end

  assign _zz_io_result_706 = _zz_io_result_701[3 : 2];
  assign _zz_io_result_707 = _zz_io_result_701[1 : 0];
  assign _zz_io_result_708 = _zz_io_result_702[3 : 2];
  assign _zz_io_result_709 = _zz_io_result_702[1 : 0];
  assign _zz_io_result_710 = (_zz_io_result_706 ^ _zz_io_result_707);
  assign _zz_io_result_711 = (_zz_io_result_708 ^ _zz_io_result_709);
  assign _zz_io_result_713 = ((_zz_io_result_711[0] && _zz_io_result_710[1]) ^ (_zz_io_result_710[0] && _zz_io_result_711[1]));
  always @(*) begin
    _zz_io_result_714[1] = ((_zz_io_result_711[0] && _zz_io_result_710[0]) ^ _zz_io_result_713);
    _zz_io_result_714[0] = ((_zz_io_result_711[1] && _zz_io_result_710[1]) ^ _zz_io_result_713);
  end

  assign _zz_io_result_712 = _zz_io_result_714;
  always @(*) begin
    _zz_io_result_716[1] = _zz_io_result_712[0];
    _zz_io_result_716[0] = (_zz_io_result_712[0] ^ _zz_io_result_712[1]);
  end

  assign _zz_io_result_715 = _zz_io_result_716;
  assign _zz_io_result_717 = ((_zz_io_result_708[0] && _zz_io_result_706[1]) ^ (_zz_io_result_706[0] && _zz_io_result_708[1]));
  always @(*) begin
    _zz_io_result_718[1] = ((_zz_io_result_708[0] && _zz_io_result_706[0]) ^ _zz_io_result_717);
    _zz_io_result_718[0] = ((_zz_io_result_708[1] && _zz_io_result_706[1]) ^ _zz_io_result_717);
  end

  assign _zz_io_result_719 = ((_zz_io_result_709[0] && _zz_io_result_707[1]) ^ (_zz_io_result_707[0] && _zz_io_result_709[1]));
  always @(*) begin
    _zz_io_result_720[1] = ((_zz_io_result_709[0] && _zz_io_result_707[0]) ^ _zz_io_result_719);
    _zz_io_result_720[0] = ((_zz_io_result_709[1] && _zz_io_result_707[1]) ^ _zz_io_result_719);
  end

  always @(*) begin
    _zz_io_result_705[3 : 2] = (_zz_io_result_718 ^ _zz_io_result_715);
    _zz_io_result_705[1 : 0] = (_zz_io_result_720 ^ _zz_io_result_715);
  end

  assign _zz_io_result_721 = (_zz_io_result_704 ^ _zz_io_result_705);
  assign _zz_io_result_724 = _zz_io_result_721[3 : 2];
  assign _zz_io_result_725 = _zz_io_result_721[1 : 0];
  assign _zz_io_result_726 = (_zz_io_result_724 ^ _zz_io_result_725);
  always @(*) begin
    _zz_io_result_727[1] = _zz_io_result_726[1];
    _zz_io_result_727[0] = (_zz_io_result_726[0] ^ _zz_io_result_726[1]);
  end

  assign _zz_io_result_728 = ((_zz_io_result_725[0] && _zz_io_result_724[1]) ^ (_zz_io_result_724[0] && _zz_io_result_725[1]));
  always @(*) begin
    _zz_io_result_729[1] = ((_zz_io_result_725[0] && _zz_io_result_724[0]) ^ _zz_io_result_728);
    _zz_io_result_729[0] = ((_zz_io_result_725[1] && _zz_io_result_724[1]) ^ _zz_io_result_728);
  end

  assign _zz_io_result_730 = (_zz_io_result_727 ^ _zz_io_result_729);
  always @(*) begin
    _zz_io_result_732[1] = _zz_io_result_730[0];
    _zz_io_result_732[0] = _zz_io_result_730[1];
  end

  assign _zz_io_result_731 = _zz_io_result_732;
  assign _zz_io_result_733 = ((_zz_io_result_731[0] && _zz_io_result_724[1]) ^ (_zz_io_result_724[0] && _zz_io_result_731[1]));
  always @(*) begin
    _zz_io_result_734[1] = ((_zz_io_result_731[0] && _zz_io_result_724[0]) ^ _zz_io_result_733);
    _zz_io_result_734[0] = ((_zz_io_result_731[1] && _zz_io_result_724[1]) ^ _zz_io_result_733);
  end

  assign _zz_io_result_735 = ((_zz_io_result_731[0] && _zz_io_result_725[1]) ^ (_zz_io_result_725[0] && _zz_io_result_731[1]));
  always @(*) begin
    _zz_io_result_736[1] = ((_zz_io_result_731[0] && _zz_io_result_725[0]) ^ _zz_io_result_735);
    _zz_io_result_736[0] = ((_zz_io_result_731[1] && _zz_io_result_725[1]) ^ _zz_io_result_735);
  end

  always @(*) begin
    _zz_io_result_723[3 : 2] = _zz_io_result_736;
    _zz_io_result_723[1 : 0] = _zz_io_result_734;
  end

  assign _zz_io_result_722 = _zz_io_result_723;
  assign _zz_io_result_738 = _zz_io_result_701[3 : 2];
  assign _zz_io_result_739 = _zz_io_result_701[1 : 0];
  assign _zz_io_result_740 = _zz_io_result_722[3 : 2];
  assign _zz_io_result_741 = _zz_io_result_722[1 : 0];
  assign _zz_io_result_742 = (_zz_io_result_738 ^ _zz_io_result_739);
  assign _zz_io_result_743 = (_zz_io_result_740 ^ _zz_io_result_741);
  assign _zz_io_result_745 = ((_zz_io_result_743[0] && _zz_io_result_742[1]) ^ (_zz_io_result_742[0] && _zz_io_result_743[1]));
  always @(*) begin
    _zz_io_result_746[1] = ((_zz_io_result_743[0] && _zz_io_result_742[0]) ^ _zz_io_result_745);
    _zz_io_result_746[0] = ((_zz_io_result_743[1] && _zz_io_result_742[1]) ^ _zz_io_result_745);
  end

  assign _zz_io_result_744 = _zz_io_result_746;
  always @(*) begin
    _zz_io_result_748[1] = _zz_io_result_744[0];
    _zz_io_result_748[0] = (_zz_io_result_744[0] ^ _zz_io_result_744[1]);
  end

  assign _zz_io_result_747 = _zz_io_result_748;
  assign _zz_io_result_749 = ((_zz_io_result_740[0] && _zz_io_result_738[1]) ^ (_zz_io_result_738[0] && _zz_io_result_740[1]));
  always @(*) begin
    _zz_io_result_750[1] = ((_zz_io_result_740[0] && _zz_io_result_738[0]) ^ _zz_io_result_749);
    _zz_io_result_750[0] = ((_zz_io_result_740[1] && _zz_io_result_738[1]) ^ _zz_io_result_749);
  end

  assign _zz_io_result_751 = ((_zz_io_result_741[0] && _zz_io_result_739[1]) ^ (_zz_io_result_739[0] && _zz_io_result_741[1]));
  always @(*) begin
    _zz_io_result_752[1] = ((_zz_io_result_741[0] && _zz_io_result_739[0]) ^ _zz_io_result_751);
    _zz_io_result_752[0] = ((_zz_io_result_741[1] && _zz_io_result_739[1]) ^ _zz_io_result_751);
  end

  always @(*) begin
    _zz_io_result_737[3 : 2] = (_zz_io_result_750 ^ _zz_io_result_747);
    _zz_io_result_737[1 : 0] = (_zz_io_result_752 ^ _zz_io_result_747);
  end

  assign _zz_io_result_754 = _zz_io_result_702[3 : 2];
  assign _zz_io_result_755 = _zz_io_result_702[1 : 0];
  assign _zz_io_result_756 = _zz_io_result_722[3 : 2];
  assign _zz_io_result_757 = _zz_io_result_722[1 : 0];
  assign _zz_io_result_758 = (_zz_io_result_754 ^ _zz_io_result_755);
  assign _zz_io_result_759 = (_zz_io_result_756 ^ _zz_io_result_757);
  assign _zz_io_result_761 = ((_zz_io_result_759[0] && _zz_io_result_758[1]) ^ (_zz_io_result_758[0] && _zz_io_result_759[1]));
  always @(*) begin
    _zz_io_result_762[1] = ((_zz_io_result_759[0] && _zz_io_result_758[0]) ^ _zz_io_result_761);
    _zz_io_result_762[0] = ((_zz_io_result_759[1] && _zz_io_result_758[1]) ^ _zz_io_result_761);
  end

  assign _zz_io_result_760 = _zz_io_result_762;
  always @(*) begin
    _zz_io_result_764[1] = _zz_io_result_760[0];
    _zz_io_result_764[0] = (_zz_io_result_760[0] ^ _zz_io_result_760[1]);
  end

  assign _zz_io_result_763 = _zz_io_result_764;
  assign _zz_io_result_765 = ((_zz_io_result_756[0] && _zz_io_result_754[1]) ^ (_zz_io_result_754[0] && _zz_io_result_756[1]));
  always @(*) begin
    _zz_io_result_766[1] = ((_zz_io_result_756[0] && _zz_io_result_754[0]) ^ _zz_io_result_765);
    _zz_io_result_766[0] = ((_zz_io_result_756[1] && _zz_io_result_754[1]) ^ _zz_io_result_765);
  end

  assign _zz_io_result_767 = ((_zz_io_result_757[0] && _zz_io_result_755[1]) ^ (_zz_io_result_755[0] && _zz_io_result_757[1]));
  always @(*) begin
    _zz_io_result_768[1] = ((_zz_io_result_757[0] && _zz_io_result_755[0]) ^ _zz_io_result_767);
    _zz_io_result_768[0] = ((_zz_io_result_757[1] && _zz_io_result_755[1]) ^ _zz_io_result_767);
  end

  always @(*) begin
    _zz_io_result_753[3 : 2] = (_zz_io_result_766 ^ _zz_io_result_763);
    _zz_io_result_753[1 : 0] = (_zz_io_result_768 ^ _zz_io_result_763);
  end

  always @(*) begin
    _zz_io_result_700[7 : 4] = _zz_io_result_753;
    _zz_io_result_700[3 : 0] = _zz_io_result_737;
  end

  assign _zz_io_result_699 = _zz_io_result_700;
  always @(*) begin
    _zz_io_result_770[7] = (_zz_io_result_699[5] ^ _zz_io_result_699[3]);
    _zz_io_result_770[6] = (_zz_io_result_699[7] ^ _zz_io_result_699[3]);
    _zz_io_result_770[5] = (_zz_io_result_699[6] ^ _zz_io_result_699[0]);
    _zz_io_result_770[4] = ((_zz_io_result_699[7] ^ _zz_io_result_699[5]) ^ _zz_io_result_699[3]);
    _zz_io_result_770[3] = ((((_zz_io_result_699[7] ^ _zz_io_result_699[6]) ^ _zz_io_result_699[5]) ^ _zz_io_result_699[4]) ^ _zz_io_result_699[3]);
    _zz_io_result_770[2] = ((((_zz_io_result_699[6] ^ _zz_io_result_699[5]) ^ _zz_io_result_699[3]) ^ _zz_io_result_699[2]) ^ _zz_io_result_699[0]);
    _zz_io_result_770[1] = ((_zz_io_result_699[5] ^ _zz_io_result_699[4]) ^ _zz_io_result_699[1]);
    _zz_io_result_770[0] = ((_zz_io_result_699[6] ^ _zz_io_result_699[4]) ^ _zz_io_result_699[1]);
  end

  assign _zz_io_result_769 = _zz_io_result_770;
  always @(*) begin
    _zz_io_result_696[7] = _zz_io_result_769[7];
    _zz_io_result_696[6] = (! _zz_io_result_769[6]);
    _zz_io_result_696[5] = (! _zz_io_result_769[5]);
    _zz_io_result_696[4] = _zz_io_result_769[4];
    _zz_io_result_696[3] = _zz_io_result_769[3];
    _zz_io_result_696[2] = _zz_io_result_769[2];
    _zz_io_result_696[1] = (! _zz_io_result_769[1]);
    _zz_io_result_696[0] = (! _zz_io_result_769[0]);
  end

  assign _zz_io_result_771 = _zz_io_result_2[23 : 16];
  always @(*) begin
    _zz_io_result_774[7] = (((((_zz_io_result_771[7] ^ _zz_io_result_771[6]) ^ _zz_io_result_771[5]) ^ _zz_io_result_771[2]) ^ _zz_io_result_771[1]) ^ _zz_io_result_771[0]);
    _zz_io_result_774[6] = (((_zz_io_result_771[6] ^ _zz_io_result_771[5]) ^ _zz_io_result_771[4]) ^ _zz_io_result_771[0]);
    _zz_io_result_774[5] = (((_zz_io_result_771[6] ^ _zz_io_result_771[5]) ^ _zz_io_result_771[1]) ^ _zz_io_result_771[0]);
    _zz_io_result_774[4] = (((_zz_io_result_771[7] ^ _zz_io_result_771[6]) ^ _zz_io_result_771[5]) ^ _zz_io_result_771[0]);
    _zz_io_result_774[3] = ((((_zz_io_result_771[7] ^ _zz_io_result_771[4]) ^ _zz_io_result_771[3]) ^ _zz_io_result_771[1]) ^ _zz_io_result_771[0]);
    _zz_io_result_774[2] = _zz_io_result_771[0];
    _zz_io_result_774[1] = ((_zz_io_result_771[6] ^ _zz_io_result_771[5]) ^ _zz_io_result_771[0]);
    _zz_io_result_774[0] = ((((_zz_io_result_771[6] ^ _zz_io_result_771[3]) ^ _zz_io_result_771[2]) ^ _zz_io_result_771[1]) ^ _zz_io_result_771[0]);
  end

  assign _zz_io_result_773 = _zz_io_result_774;
  assign _zz_io_result_777 = _zz_io_result_773[7 : 4];
  assign _zz_io_result_778 = _zz_io_result_773[3 : 0];
  assign _zz_io_result_779 = (_zz_io_result_777 ^ _zz_io_result_778);
  always @(*) begin
    _zz_io_result_780[3] = (_zz_io_result_779[2] ^ _zz_io_result_779[0]);
    _zz_io_result_780[2] = (_zz_io_result_779[3] ^ _zz_io_result_779[1]);
    _zz_io_result_780[1] = (_zz_io_result_779[1] ^ _zz_io_result_779[0]);
    _zz_io_result_780[0] = _zz_io_result_779[0];
  end

  assign _zz_io_result_782 = _zz_io_result_777[3 : 2];
  assign _zz_io_result_783 = _zz_io_result_777[1 : 0];
  assign _zz_io_result_784 = _zz_io_result_778[3 : 2];
  assign _zz_io_result_785 = _zz_io_result_778[1 : 0];
  assign _zz_io_result_786 = (_zz_io_result_782 ^ _zz_io_result_783);
  assign _zz_io_result_787 = (_zz_io_result_784 ^ _zz_io_result_785);
  assign _zz_io_result_789 = ((_zz_io_result_787[0] && _zz_io_result_786[1]) ^ (_zz_io_result_786[0] && _zz_io_result_787[1]));
  always @(*) begin
    _zz_io_result_790[1] = ((_zz_io_result_787[0] && _zz_io_result_786[0]) ^ _zz_io_result_789);
    _zz_io_result_790[0] = ((_zz_io_result_787[1] && _zz_io_result_786[1]) ^ _zz_io_result_789);
  end

  assign _zz_io_result_788 = _zz_io_result_790;
  always @(*) begin
    _zz_io_result_792[1] = _zz_io_result_788[0];
    _zz_io_result_792[0] = (_zz_io_result_788[0] ^ _zz_io_result_788[1]);
  end

  assign _zz_io_result_791 = _zz_io_result_792;
  assign _zz_io_result_793 = ((_zz_io_result_784[0] && _zz_io_result_782[1]) ^ (_zz_io_result_782[0] && _zz_io_result_784[1]));
  always @(*) begin
    _zz_io_result_794[1] = ((_zz_io_result_784[0] && _zz_io_result_782[0]) ^ _zz_io_result_793);
    _zz_io_result_794[0] = ((_zz_io_result_784[1] && _zz_io_result_782[1]) ^ _zz_io_result_793);
  end

  assign _zz_io_result_795 = ((_zz_io_result_785[0] && _zz_io_result_783[1]) ^ (_zz_io_result_783[0] && _zz_io_result_785[1]));
  always @(*) begin
    _zz_io_result_796[1] = ((_zz_io_result_785[0] && _zz_io_result_783[0]) ^ _zz_io_result_795);
    _zz_io_result_796[0] = ((_zz_io_result_785[1] && _zz_io_result_783[1]) ^ _zz_io_result_795);
  end

  always @(*) begin
    _zz_io_result_781[3 : 2] = (_zz_io_result_794 ^ _zz_io_result_791);
    _zz_io_result_781[1 : 0] = (_zz_io_result_796 ^ _zz_io_result_791);
  end

  assign _zz_io_result_797 = (_zz_io_result_780 ^ _zz_io_result_781);
  assign _zz_io_result_800 = _zz_io_result_797[3 : 2];
  assign _zz_io_result_801 = _zz_io_result_797[1 : 0];
  assign _zz_io_result_802 = (_zz_io_result_800 ^ _zz_io_result_801);
  always @(*) begin
    _zz_io_result_803[1] = _zz_io_result_802[1];
    _zz_io_result_803[0] = (_zz_io_result_802[0] ^ _zz_io_result_802[1]);
  end

  assign _zz_io_result_804 = ((_zz_io_result_801[0] && _zz_io_result_800[1]) ^ (_zz_io_result_800[0] && _zz_io_result_801[1]));
  always @(*) begin
    _zz_io_result_805[1] = ((_zz_io_result_801[0] && _zz_io_result_800[0]) ^ _zz_io_result_804);
    _zz_io_result_805[0] = ((_zz_io_result_801[1] && _zz_io_result_800[1]) ^ _zz_io_result_804);
  end

  assign _zz_io_result_806 = (_zz_io_result_803 ^ _zz_io_result_805);
  always @(*) begin
    _zz_io_result_808[1] = _zz_io_result_806[0];
    _zz_io_result_808[0] = _zz_io_result_806[1];
  end

  assign _zz_io_result_807 = _zz_io_result_808;
  assign _zz_io_result_809 = ((_zz_io_result_807[0] && _zz_io_result_800[1]) ^ (_zz_io_result_800[0] && _zz_io_result_807[1]));
  always @(*) begin
    _zz_io_result_810[1] = ((_zz_io_result_807[0] && _zz_io_result_800[0]) ^ _zz_io_result_809);
    _zz_io_result_810[0] = ((_zz_io_result_807[1] && _zz_io_result_800[1]) ^ _zz_io_result_809);
  end

  assign _zz_io_result_811 = ((_zz_io_result_807[0] && _zz_io_result_801[1]) ^ (_zz_io_result_801[0] && _zz_io_result_807[1]));
  always @(*) begin
    _zz_io_result_812[1] = ((_zz_io_result_807[0] && _zz_io_result_801[0]) ^ _zz_io_result_811);
    _zz_io_result_812[0] = ((_zz_io_result_807[1] && _zz_io_result_801[1]) ^ _zz_io_result_811);
  end

  always @(*) begin
    _zz_io_result_799[3 : 2] = _zz_io_result_812;
    _zz_io_result_799[1 : 0] = _zz_io_result_810;
  end

  assign _zz_io_result_798 = _zz_io_result_799;
  assign _zz_io_result_814 = _zz_io_result_777[3 : 2];
  assign _zz_io_result_815 = _zz_io_result_777[1 : 0];
  assign _zz_io_result_816 = _zz_io_result_798[3 : 2];
  assign _zz_io_result_817 = _zz_io_result_798[1 : 0];
  assign _zz_io_result_818 = (_zz_io_result_814 ^ _zz_io_result_815);
  assign _zz_io_result_819 = (_zz_io_result_816 ^ _zz_io_result_817);
  assign _zz_io_result_821 = ((_zz_io_result_819[0] && _zz_io_result_818[1]) ^ (_zz_io_result_818[0] && _zz_io_result_819[1]));
  always @(*) begin
    _zz_io_result_822[1] = ((_zz_io_result_819[0] && _zz_io_result_818[0]) ^ _zz_io_result_821);
    _zz_io_result_822[0] = ((_zz_io_result_819[1] && _zz_io_result_818[1]) ^ _zz_io_result_821);
  end

  assign _zz_io_result_820 = _zz_io_result_822;
  always @(*) begin
    _zz_io_result_824[1] = _zz_io_result_820[0];
    _zz_io_result_824[0] = (_zz_io_result_820[0] ^ _zz_io_result_820[1]);
  end

  assign _zz_io_result_823 = _zz_io_result_824;
  assign _zz_io_result_825 = ((_zz_io_result_816[0] && _zz_io_result_814[1]) ^ (_zz_io_result_814[0] && _zz_io_result_816[1]));
  always @(*) begin
    _zz_io_result_826[1] = ((_zz_io_result_816[0] && _zz_io_result_814[0]) ^ _zz_io_result_825);
    _zz_io_result_826[0] = ((_zz_io_result_816[1] && _zz_io_result_814[1]) ^ _zz_io_result_825);
  end

  assign _zz_io_result_827 = ((_zz_io_result_817[0] && _zz_io_result_815[1]) ^ (_zz_io_result_815[0] && _zz_io_result_817[1]));
  always @(*) begin
    _zz_io_result_828[1] = ((_zz_io_result_817[0] && _zz_io_result_815[0]) ^ _zz_io_result_827);
    _zz_io_result_828[0] = ((_zz_io_result_817[1] && _zz_io_result_815[1]) ^ _zz_io_result_827);
  end

  always @(*) begin
    _zz_io_result_813[3 : 2] = (_zz_io_result_826 ^ _zz_io_result_823);
    _zz_io_result_813[1 : 0] = (_zz_io_result_828 ^ _zz_io_result_823);
  end

  assign _zz_io_result_830 = _zz_io_result_778[3 : 2];
  assign _zz_io_result_831 = _zz_io_result_778[1 : 0];
  assign _zz_io_result_832 = _zz_io_result_798[3 : 2];
  assign _zz_io_result_833 = _zz_io_result_798[1 : 0];
  assign _zz_io_result_834 = (_zz_io_result_830 ^ _zz_io_result_831);
  assign _zz_io_result_835 = (_zz_io_result_832 ^ _zz_io_result_833);
  assign _zz_io_result_837 = ((_zz_io_result_835[0] && _zz_io_result_834[1]) ^ (_zz_io_result_834[0] && _zz_io_result_835[1]));
  always @(*) begin
    _zz_io_result_838[1] = ((_zz_io_result_835[0] && _zz_io_result_834[0]) ^ _zz_io_result_837);
    _zz_io_result_838[0] = ((_zz_io_result_835[1] && _zz_io_result_834[1]) ^ _zz_io_result_837);
  end

  assign _zz_io_result_836 = _zz_io_result_838;
  always @(*) begin
    _zz_io_result_840[1] = _zz_io_result_836[0];
    _zz_io_result_840[0] = (_zz_io_result_836[0] ^ _zz_io_result_836[1]);
  end

  assign _zz_io_result_839 = _zz_io_result_840;
  assign _zz_io_result_841 = ((_zz_io_result_832[0] && _zz_io_result_830[1]) ^ (_zz_io_result_830[0] && _zz_io_result_832[1]));
  always @(*) begin
    _zz_io_result_842[1] = ((_zz_io_result_832[0] && _zz_io_result_830[0]) ^ _zz_io_result_841);
    _zz_io_result_842[0] = ((_zz_io_result_832[1] && _zz_io_result_830[1]) ^ _zz_io_result_841);
  end

  assign _zz_io_result_843 = ((_zz_io_result_833[0] && _zz_io_result_831[1]) ^ (_zz_io_result_831[0] && _zz_io_result_833[1]));
  always @(*) begin
    _zz_io_result_844[1] = ((_zz_io_result_833[0] && _zz_io_result_831[0]) ^ _zz_io_result_843);
    _zz_io_result_844[0] = ((_zz_io_result_833[1] && _zz_io_result_831[1]) ^ _zz_io_result_843);
  end

  always @(*) begin
    _zz_io_result_829[3 : 2] = (_zz_io_result_842 ^ _zz_io_result_839);
    _zz_io_result_829[1 : 0] = (_zz_io_result_844 ^ _zz_io_result_839);
  end

  always @(*) begin
    _zz_io_result_776[7 : 4] = _zz_io_result_829;
    _zz_io_result_776[3 : 0] = _zz_io_result_813;
  end

  assign _zz_io_result_775 = _zz_io_result_776;
  always @(*) begin
    _zz_io_result_846[7] = (_zz_io_result_775[5] ^ _zz_io_result_775[3]);
    _zz_io_result_846[6] = (_zz_io_result_775[7] ^ _zz_io_result_775[3]);
    _zz_io_result_846[5] = (_zz_io_result_775[6] ^ _zz_io_result_775[0]);
    _zz_io_result_846[4] = ((_zz_io_result_775[7] ^ _zz_io_result_775[5]) ^ _zz_io_result_775[3]);
    _zz_io_result_846[3] = ((((_zz_io_result_775[7] ^ _zz_io_result_775[6]) ^ _zz_io_result_775[5]) ^ _zz_io_result_775[4]) ^ _zz_io_result_775[3]);
    _zz_io_result_846[2] = ((((_zz_io_result_775[6] ^ _zz_io_result_775[5]) ^ _zz_io_result_775[3]) ^ _zz_io_result_775[2]) ^ _zz_io_result_775[0]);
    _zz_io_result_846[1] = ((_zz_io_result_775[5] ^ _zz_io_result_775[4]) ^ _zz_io_result_775[1]);
    _zz_io_result_846[0] = ((_zz_io_result_775[6] ^ _zz_io_result_775[4]) ^ _zz_io_result_775[1]);
  end

  assign _zz_io_result_845 = _zz_io_result_846;
  always @(*) begin
    _zz_io_result_772[7] = _zz_io_result_845[7];
    _zz_io_result_772[6] = (! _zz_io_result_845[6]);
    _zz_io_result_772[5] = (! _zz_io_result_845[5]);
    _zz_io_result_772[4] = _zz_io_result_845[4];
    _zz_io_result_772[3] = _zz_io_result_845[3];
    _zz_io_result_772[2] = _zz_io_result_845[2];
    _zz_io_result_772[1] = (! _zz_io_result_845[1]);
    _zz_io_result_772[0] = (! _zz_io_result_845[0]);
  end

  assign _zz_io_result_847 = _zz_io_result_2[31 : 24];
  always @(*) begin
    _zz_io_result_850[7] = (((((_zz_io_result_847[7] ^ _zz_io_result_847[6]) ^ _zz_io_result_847[5]) ^ _zz_io_result_847[2]) ^ _zz_io_result_847[1]) ^ _zz_io_result_847[0]);
    _zz_io_result_850[6] = (((_zz_io_result_847[6] ^ _zz_io_result_847[5]) ^ _zz_io_result_847[4]) ^ _zz_io_result_847[0]);
    _zz_io_result_850[5] = (((_zz_io_result_847[6] ^ _zz_io_result_847[5]) ^ _zz_io_result_847[1]) ^ _zz_io_result_847[0]);
    _zz_io_result_850[4] = (((_zz_io_result_847[7] ^ _zz_io_result_847[6]) ^ _zz_io_result_847[5]) ^ _zz_io_result_847[0]);
    _zz_io_result_850[3] = ((((_zz_io_result_847[7] ^ _zz_io_result_847[4]) ^ _zz_io_result_847[3]) ^ _zz_io_result_847[1]) ^ _zz_io_result_847[0]);
    _zz_io_result_850[2] = _zz_io_result_847[0];
    _zz_io_result_850[1] = ((_zz_io_result_847[6] ^ _zz_io_result_847[5]) ^ _zz_io_result_847[0]);
    _zz_io_result_850[0] = ((((_zz_io_result_847[6] ^ _zz_io_result_847[3]) ^ _zz_io_result_847[2]) ^ _zz_io_result_847[1]) ^ _zz_io_result_847[0]);
  end

  assign _zz_io_result_849 = _zz_io_result_850;
  assign _zz_io_result_853 = _zz_io_result_849[7 : 4];
  assign _zz_io_result_854 = _zz_io_result_849[3 : 0];
  assign _zz_io_result_855 = (_zz_io_result_853 ^ _zz_io_result_854);
  always @(*) begin
    _zz_io_result_856[3] = (_zz_io_result_855[2] ^ _zz_io_result_855[0]);
    _zz_io_result_856[2] = (_zz_io_result_855[3] ^ _zz_io_result_855[1]);
    _zz_io_result_856[1] = (_zz_io_result_855[1] ^ _zz_io_result_855[0]);
    _zz_io_result_856[0] = _zz_io_result_855[0];
  end

  assign _zz_io_result_858 = _zz_io_result_853[3 : 2];
  assign _zz_io_result_859 = _zz_io_result_853[1 : 0];
  assign _zz_io_result_860 = _zz_io_result_854[3 : 2];
  assign _zz_io_result_861 = _zz_io_result_854[1 : 0];
  assign _zz_io_result_862 = (_zz_io_result_858 ^ _zz_io_result_859);
  assign _zz_io_result_863 = (_zz_io_result_860 ^ _zz_io_result_861);
  assign _zz_io_result_865 = ((_zz_io_result_863[0] && _zz_io_result_862[1]) ^ (_zz_io_result_862[0] && _zz_io_result_863[1]));
  always @(*) begin
    _zz_io_result_866[1] = ((_zz_io_result_863[0] && _zz_io_result_862[0]) ^ _zz_io_result_865);
    _zz_io_result_866[0] = ((_zz_io_result_863[1] && _zz_io_result_862[1]) ^ _zz_io_result_865);
  end

  assign _zz_io_result_864 = _zz_io_result_866;
  always @(*) begin
    _zz_io_result_868[1] = _zz_io_result_864[0];
    _zz_io_result_868[0] = (_zz_io_result_864[0] ^ _zz_io_result_864[1]);
  end

  assign _zz_io_result_867 = _zz_io_result_868;
  assign _zz_io_result_869 = ((_zz_io_result_860[0] && _zz_io_result_858[1]) ^ (_zz_io_result_858[0] && _zz_io_result_860[1]));
  always @(*) begin
    _zz_io_result_870[1] = ((_zz_io_result_860[0] && _zz_io_result_858[0]) ^ _zz_io_result_869);
    _zz_io_result_870[0] = ((_zz_io_result_860[1] && _zz_io_result_858[1]) ^ _zz_io_result_869);
  end

  assign _zz_io_result_871 = ((_zz_io_result_861[0] && _zz_io_result_859[1]) ^ (_zz_io_result_859[0] && _zz_io_result_861[1]));
  always @(*) begin
    _zz_io_result_872[1] = ((_zz_io_result_861[0] && _zz_io_result_859[0]) ^ _zz_io_result_871);
    _zz_io_result_872[0] = ((_zz_io_result_861[1] && _zz_io_result_859[1]) ^ _zz_io_result_871);
  end

  always @(*) begin
    _zz_io_result_857[3 : 2] = (_zz_io_result_870 ^ _zz_io_result_867);
    _zz_io_result_857[1 : 0] = (_zz_io_result_872 ^ _zz_io_result_867);
  end

  assign _zz_io_result_873 = (_zz_io_result_856 ^ _zz_io_result_857);
  assign _zz_io_result_876 = _zz_io_result_873[3 : 2];
  assign _zz_io_result_877 = _zz_io_result_873[1 : 0];
  assign _zz_io_result_878 = (_zz_io_result_876 ^ _zz_io_result_877);
  always @(*) begin
    _zz_io_result_879[1] = _zz_io_result_878[1];
    _zz_io_result_879[0] = (_zz_io_result_878[0] ^ _zz_io_result_878[1]);
  end

  assign _zz_io_result_880 = ((_zz_io_result_877[0] && _zz_io_result_876[1]) ^ (_zz_io_result_876[0] && _zz_io_result_877[1]));
  always @(*) begin
    _zz_io_result_881[1] = ((_zz_io_result_877[0] && _zz_io_result_876[0]) ^ _zz_io_result_880);
    _zz_io_result_881[0] = ((_zz_io_result_877[1] && _zz_io_result_876[1]) ^ _zz_io_result_880);
  end

  assign _zz_io_result_882 = (_zz_io_result_879 ^ _zz_io_result_881);
  always @(*) begin
    _zz_io_result_884[1] = _zz_io_result_882[0];
    _zz_io_result_884[0] = _zz_io_result_882[1];
  end

  assign _zz_io_result_883 = _zz_io_result_884;
  assign _zz_io_result_885 = ((_zz_io_result_883[0] && _zz_io_result_876[1]) ^ (_zz_io_result_876[0] && _zz_io_result_883[1]));
  always @(*) begin
    _zz_io_result_886[1] = ((_zz_io_result_883[0] && _zz_io_result_876[0]) ^ _zz_io_result_885);
    _zz_io_result_886[0] = ((_zz_io_result_883[1] && _zz_io_result_876[1]) ^ _zz_io_result_885);
  end

  assign _zz_io_result_887 = ((_zz_io_result_883[0] && _zz_io_result_877[1]) ^ (_zz_io_result_877[0] && _zz_io_result_883[1]));
  always @(*) begin
    _zz_io_result_888[1] = ((_zz_io_result_883[0] && _zz_io_result_877[0]) ^ _zz_io_result_887);
    _zz_io_result_888[0] = ((_zz_io_result_883[1] && _zz_io_result_877[1]) ^ _zz_io_result_887);
  end

  always @(*) begin
    _zz_io_result_875[3 : 2] = _zz_io_result_888;
    _zz_io_result_875[1 : 0] = _zz_io_result_886;
  end

  assign _zz_io_result_874 = _zz_io_result_875;
  assign _zz_io_result_890 = _zz_io_result_853[3 : 2];
  assign _zz_io_result_891 = _zz_io_result_853[1 : 0];
  assign _zz_io_result_892 = _zz_io_result_874[3 : 2];
  assign _zz_io_result_893 = _zz_io_result_874[1 : 0];
  assign _zz_io_result_894 = (_zz_io_result_890 ^ _zz_io_result_891);
  assign _zz_io_result_895 = (_zz_io_result_892 ^ _zz_io_result_893);
  assign _zz_io_result_897 = ((_zz_io_result_895[0] && _zz_io_result_894[1]) ^ (_zz_io_result_894[0] && _zz_io_result_895[1]));
  always @(*) begin
    _zz_io_result_898[1] = ((_zz_io_result_895[0] && _zz_io_result_894[0]) ^ _zz_io_result_897);
    _zz_io_result_898[0] = ((_zz_io_result_895[1] && _zz_io_result_894[1]) ^ _zz_io_result_897);
  end

  assign _zz_io_result_896 = _zz_io_result_898;
  always @(*) begin
    _zz_io_result_900[1] = _zz_io_result_896[0];
    _zz_io_result_900[0] = (_zz_io_result_896[0] ^ _zz_io_result_896[1]);
  end

  assign _zz_io_result_899 = _zz_io_result_900;
  assign _zz_io_result_901 = ((_zz_io_result_892[0] && _zz_io_result_890[1]) ^ (_zz_io_result_890[0] && _zz_io_result_892[1]));
  always @(*) begin
    _zz_io_result_902[1] = ((_zz_io_result_892[0] && _zz_io_result_890[0]) ^ _zz_io_result_901);
    _zz_io_result_902[0] = ((_zz_io_result_892[1] && _zz_io_result_890[1]) ^ _zz_io_result_901);
  end

  assign _zz_io_result_903 = ((_zz_io_result_893[0] && _zz_io_result_891[1]) ^ (_zz_io_result_891[0] && _zz_io_result_893[1]));
  always @(*) begin
    _zz_io_result_904[1] = ((_zz_io_result_893[0] && _zz_io_result_891[0]) ^ _zz_io_result_903);
    _zz_io_result_904[0] = ((_zz_io_result_893[1] && _zz_io_result_891[1]) ^ _zz_io_result_903);
  end

  always @(*) begin
    _zz_io_result_889[3 : 2] = (_zz_io_result_902 ^ _zz_io_result_899);
    _zz_io_result_889[1 : 0] = (_zz_io_result_904 ^ _zz_io_result_899);
  end

  assign _zz_io_result_906 = _zz_io_result_854[3 : 2];
  assign _zz_io_result_907 = _zz_io_result_854[1 : 0];
  assign _zz_io_result_908 = _zz_io_result_874[3 : 2];
  assign _zz_io_result_909 = _zz_io_result_874[1 : 0];
  assign _zz_io_result_910 = (_zz_io_result_906 ^ _zz_io_result_907);
  assign _zz_io_result_911 = (_zz_io_result_908 ^ _zz_io_result_909);
  assign _zz_io_result_913 = ((_zz_io_result_911[0] && _zz_io_result_910[1]) ^ (_zz_io_result_910[0] && _zz_io_result_911[1]));
  always @(*) begin
    _zz_io_result_914[1] = ((_zz_io_result_911[0] && _zz_io_result_910[0]) ^ _zz_io_result_913);
    _zz_io_result_914[0] = ((_zz_io_result_911[1] && _zz_io_result_910[1]) ^ _zz_io_result_913);
  end

  assign _zz_io_result_912 = _zz_io_result_914;
  always @(*) begin
    _zz_io_result_916[1] = _zz_io_result_912[0];
    _zz_io_result_916[0] = (_zz_io_result_912[0] ^ _zz_io_result_912[1]);
  end

  assign _zz_io_result_915 = _zz_io_result_916;
  assign _zz_io_result_917 = ((_zz_io_result_908[0] && _zz_io_result_906[1]) ^ (_zz_io_result_906[0] && _zz_io_result_908[1]));
  always @(*) begin
    _zz_io_result_918[1] = ((_zz_io_result_908[0] && _zz_io_result_906[0]) ^ _zz_io_result_917);
    _zz_io_result_918[0] = ((_zz_io_result_908[1] && _zz_io_result_906[1]) ^ _zz_io_result_917);
  end

  assign _zz_io_result_919 = ((_zz_io_result_909[0] && _zz_io_result_907[1]) ^ (_zz_io_result_907[0] && _zz_io_result_909[1]));
  always @(*) begin
    _zz_io_result_920[1] = ((_zz_io_result_909[0] && _zz_io_result_907[0]) ^ _zz_io_result_919);
    _zz_io_result_920[0] = ((_zz_io_result_909[1] && _zz_io_result_907[1]) ^ _zz_io_result_919);
  end

  always @(*) begin
    _zz_io_result_905[3 : 2] = (_zz_io_result_918 ^ _zz_io_result_915);
    _zz_io_result_905[1 : 0] = (_zz_io_result_920 ^ _zz_io_result_915);
  end

  always @(*) begin
    _zz_io_result_852[7 : 4] = _zz_io_result_905;
    _zz_io_result_852[3 : 0] = _zz_io_result_889;
  end

  assign _zz_io_result_851 = _zz_io_result_852;
  always @(*) begin
    _zz_io_result_922[7] = (_zz_io_result_851[5] ^ _zz_io_result_851[3]);
    _zz_io_result_922[6] = (_zz_io_result_851[7] ^ _zz_io_result_851[3]);
    _zz_io_result_922[5] = (_zz_io_result_851[6] ^ _zz_io_result_851[0]);
    _zz_io_result_922[4] = ((_zz_io_result_851[7] ^ _zz_io_result_851[5]) ^ _zz_io_result_851[3]);
    _zz_io_result_922[3] = ((((_zz_io_result_851[7] ^ _zz_io_result_851[6]) ^ _zz_io_result_851[5]) ^ _zz_io_result_851[4]) ^ _zz_io_result_851[3]);
    _zz_io_result_922[2] = ((((_zz_io_result_851[6] ^ _zz_io_result_851[5]) ^ _zz_io_result_851[3]) ^ _zz_io_result_851[2]) ^ _zz_io_result_851[0]);
    _zz_io_result_922[1] = ((_zz_io_result_851[5] ^ _zz_io_result_851[4]) ^ _zz_io_result_851[1]);
    _zz_io_result_922[0] = ((_zz_io_result_851[6] ^ _zz_io_result_851[4]) ^ _zz_io_result_851[1]);
  end

  assign _zz_io_result_921 = _zz_io_result_922;
  always @(*) begin
    _zz_io_result_848[7] = _zz_io_result_921[7];
    _zz_io_result_848[6] = (! _zz_io_result_921[6]);
    _zz_io_result_848[5] = (! _zz_io_result_921[5]);
    _zz_io_result_848[4] = _zz_io_result_921[4];
    _zz_io_result_848[3] = _zz_io_result_921[3];
    _zz_io_result_848[2] = _zz_io_result_921[2];
    _zz_io_result_848[1] = (! _zz_io_result_921[1]);
    _zz_io_result_848[0] = (! _zz_io_result_921[0]);
  end

  assign _zz_io_result_924 = _zz_io_result_3[7 : 0];
  always @(*) begin
    _zz_io_result_927[7] = (((((_zz_io_result_924[7] ^ _zz_io_result_924[6]) ^ _zz_io_result_924[5]) ^ _zz_io_result_924[2]) ^ _zz_io_result_924[1]) ^ _zz_io_result_924[0]);
    _zz_io_result_927[6] = (((_zz_io_result_924[6] ^ _zz_io_result_924[5]) ^ _zz_io_result_924[4]) ^ _zz_io_result_924[0]);
    _zz_io_result_927[5] = (((_zz_io_result_924[6] ^ _zz_io_result_924[5]) ^ _zz_io_result_924[1]) ^ _zz_io_result_924[0]);
    _zz_io_result_927[4] = (((_zz_io_result_924[7] ^ _zz_io_result_924[6]) ^ _zz_io_result_924[5]) ^ _zz_io_result_924[0]);
    _zz_io_result_927[3] = ((((_zz_io_result_924[7] ^ _zz_io_result_924[4]) ^ _zz_io_result_924[3]) ^ _zz_io_result_924[1]) ^ _zz_io_result_924[0]);
    _zz_io_result_927[2] = _zz_io_result_924[0];
    _zz_io_result_927[1] = ((_zz_io_result_924[6] ^ _zz_io_result_924[5]) ^ _zz_io_result_924[0]);
    _zz_io_result_927[0] = ((((_zz_io_result_924[6] ^ _zz_io_result_924[3]) ^ _zz_io_result_924[2]) ^ _zz_io_result_924[1]) ^ _zz_io_result_924[0]);
  end

  assign _zz_io_result_926 = _zz_io_result_927;
  assign _zz_io_result_930 = _zz_io_result_926[7 : 4];
  assign _zz_io_result_931 = _zz_io_result_926[3 : 0];
  assign _zz_io_result_932 = (_zz_io_result_930 ^ _zz_io_result_931);
  always @(*) begin
    _zz_io_result_933[3] = (_zz_io_result_932[2] ^ _zz_io_result_932[0]);
    _zz_io_result_933[2] = (_zz_io_result_932[3] ^ _zz_io_result_932[1]);
    _zz_io_result_933[1] = (_zz_io_result_932[1] ^ _zz_io_result_932[0]);
    _zz_io_result_933[0] = _zz_io_result_932[0];
  end

  assign _zz_io_result_935 = _zz_io_result_930[3 : 2];
  assign _zz_io_result_936 = _zz_io_result_930[1 : 0];
  assign _zz_io_result_937 = _zz_io_result_931[3 : 2];
  assign _zz_io_result_938 = _zz_io_result_931[1 : 0];
  assign _zz_io_result_939 = (_zz_io_result_935 ^ _zz_io_result_936);
  assign _zz_io_result_940 = (_zz_io_result_937 ^ _zz_io_result_938);
  assign _zz_io_result_942 = ((_zz_io_result_940[0] && _zz_io_result_939[1]) ^ (_zz_io_result_939[0] && _zz_io_result_940[1]));
  always @(*) begin
    _zz_io_result_943[1] = ((_zz_io_result_940[0] && _zz_io_result_939[0]) ^ _zz_io_result_942);
    _zz_io_result_943[0] = ((_zz_io_result_940[1] && _zz_io_result_939[1]) ^ _zz_io_result_942);
  end

  assign _zz_io_result_941 = _zz_io_result_943;
  always @(*) begin
    _zz_io_result_945[1] = _zz_io_result_941[0];
    _zz_io_result_945[0] = (_zz_io_result_941[0] ^ _zz_io_result_941[1]);
  end

  assign _zz_io_result_944 = _zz_io_result_945;
  assign _zz_io_result_946 = ((_zz_io_result_937[0] && _zz_io_result_935[1]) ^ (_zz_io_result_935[0] && _zz_io_result_937[1]));
  always @(*) begin
    _zz_io_result_947[1] = ((_zz_io_result_937[0] && _zz_io_result_935[0]) ^ _zz_io_result_946);
    _zz_io_result_947[0] = ((_zz_io_result_937[1] && _zz_io_result_935[1]) ^ _zz_io_result_946);
  end

  assign _zz_io_result_948 = ((_zz_io_result_938[0] && _zz_io_result_936[1]) ^ (_zz_io_result_936[0] && _zz_io_result_938[1]));
  always @(*) begin
    _zz_io_result_949[1] = ((_zz_io_result_938[0] && _zz_io_result_936[0]) ^ _zz_io_result_948);
    _zz_io_result_949[0] = ((_zz_io_result_938[1] && _zz_io_result_936[1]) ^ _zz_io_result_948);
  end

  always @(*) begin
    _zz_io_result_934[3 : 2] = (_zz_io_result_947 ^ _zz_io_result_944);
    _zz_io_result_934[1 : 0] = (_zz_io_result_949 ^ _zz_io_result_944);
  end

  assign _zz_io_result_950 = (_zz_io_result_933 ^ _zz_io_result_934);
  assign _zz_io_result_953 = _zz_io_result_950[3 : 2];
  assign _zz_io_result_954 = _zz_io_result_950[1 : 0];
  assign _zz_io_result_955 = (_zz_io_result_953 ^ _zz_io_result_954);
  always @(*) begin
    _zz_io_result_956[1] = _zz_io_result_955[1];
    _zz_io_result_956[0] = (_zz_io_result_955[0] ^ _zz_io_result_955[1]);
  end

  assign _zz_io_result_957 = ((_zz_io_result_954[0] && _zz_io_result_953[1]) ^ (_zz_io_result_953[0] && _zz_io_result_954[1]));
  always @(*) begin
    _zz_io_result_958[1] = ((_zz_io_result_954[0] && _zz_io_result_953[0]) ^ _zz_io_result_957);
    _zz_io_result_958[0] = ((_zz_io_result_954[1] && _zz_io_result_953[1]) ^ _zz_io_result_957);
  end

  assign _zz_io_result_959 = (_zz_io_result_956 ^ _zz_io_result_958);
  always @(*) begin
    _zz_io_result_961[1] = _zz_io_result_959[0];
    _zz_io_result_961[0] = _zz_io_result_959[1];
  end

  assign _zz_io_result_960 = _zz_io_result_961;
  assign _zz_io_result_962 = ((_zz_io_result_960[0] && _zz_io_result_953[1]) ^ (_zz_io_result_953[0] && _zz_io_result_960[1]));
  always @(*) begin
    _zz_io_result_963[1] = ((_zz_io_result_960[0] && _zz_io_result_953[0]) ^ _zz_io_result_962);
    _zz_io_result_963[0] = ((_zz_io_result_960[1] && _zz_io_result_953[1]) ^ _zz_io_result_962);
  end

  assign _zz_io_result_964 = ((_zz_io_result_960[0] && _zz_io_result_954[1]) ^ (_zz_io_result_954[0] && _zz_io_result_960[1]));
  always @(*) begin
    _zz_io_result_965[1] = ((_zz_io_result_960[0] && _zz_io_result_954[0]) ^ _zz_io_result_964);
    _zz_io_result_965[0] = ((_zz_io_result_960[1] && _zz_io_result_954[1]) ^ _zz_io_result_964);
  end

  always @(*) begin
    _zz_io_result_952[3 : 2] = _zz_io_result_965;
    _zz_io_result_952[1 : 0] = _zz_io_result_963;
  end

  assign _zz_io_result_951 = _zz_io_result_952;
  assign _zz_io_result_967 = _zz_io_result_930[3 : 2];
  assign _zz_io_result_968 = _zz_io_result_930[1 : 0];
  assign _zz_io_result_969 = _zz_io_result_951[3 : 2];
  assign _zz_io_result_970 = _zz_io_result_951[1 : 0];
  assign _zz_io_result_971 = (_zz_io_result_967 ^ _zz_io_result_968);
  assign _zz_io_result_972 = (_zz_io_result_969 ^ _zz_io_result_970);
  assign _zz_io_result_974 = ((_zz_io_result_972[0] && _zz_io_result_971[1]) ^ (_zz_io_result_971[0] && _zz_io_result_972[1]));
  always @(*) begin
    _zz_io_result_975[1] = ((_zz_io_result_972[0] && _zz_io_result_971[0]) ^ _zz_io_result_974);
    _zz_io_result_975[0] = ((_zz_io_result_972[1] && _zz_io_result_971[1]) ^ _zz_io_result_974);
  end

  assign _zz_io_result_973 = _zz_io_result_975;
  always @(*) begin
    _zz_io_result_977[1] = _zz_io_result_973[0];
    _zz_io_result_977[0] = (_zz_io_result_973[0] ^ _zz_io_result_973[1]);
  end

  assign _zz_io_result_976 = _zz_io_result_977;
  assign _zz_io_result_978 = ((_zz_io_result_969[0] && _zz_io_result_967[1]) ^ (_zz_io_result_967[0] && _zz_io_result_969[1]));
  always @(*) begin
    _zz_io_result_979[1] = ((_zz_io_result_969[0] && _zz_io_result_967[0]) ^ _zz_io_result_978);
    _zz_io_result_979[0] = ((_zz_io_result_969[1] && _zz_io_result_967[1]) ^ _zz_io_result_978);
  end

  assign _zz_io_result_980 = ((_zz_io_result_970[0] && _zz_io_result_968[1]) ^ (_zz_io_result_968[0] && _zz_io_result_970[1]));
  always @(*) begin
    _zz_io_result_981[1] = ((_zz_io_result_970[0] && _zz_io_result_968[0]) ^ _zz_io_result_980);
    _zz_io_result_981[0] = ((_zz_io_result_970[1] && _zz_io_result_968[1]) ^ _zz_io_result_980);
  end

  always @(*) begin
    _zz_io_result_966[3 : 2] = (_zz_io_result_979 ^ _zz_io_result_976);
    _zz_io_result_966[1 : 0] = (_zz_io_result_981 ^ _zz_io_result_976);
  end

  assign _zz_io_result_983 = _zz_io_result_931[3 : 2];
  assign _zz_io_result_984 = _zz_io_result_931[1 : 0];
  assign _zz_io_result_985 = _zz_io_result_951[3 : 2];
  assign _zz_io_result_986 = _zz_io_result_951[1 : 0];
  assign _zz_io_result_987 = (_zz_io_result_983 ^ _zz_io_result_984);
  assign _zz_io_result_988 = (_zz_io_result_985 ^ _zz_io_result_986);
  assign _zz_io_result_990 = ((_zz_io_result_988[0] && _zz_io_result_987[1]) ^ (_zz_io_result_987[0] && _zz_io_result_988[1]));
  always @(*) begin
    _zz_io_result_991[1] = ((_zz_io_result_988[0] && _zz_io_result_987[0]) ^ _zz_io_result_990);
    _zz_io_result_991[0] = ((_zz_io_result_988[1] && _zz_io_result_987[1]) ^ _zz_io_result_990);
  end

  assign _zz_io_result_989 = _zz_io_result_991;
  always @(*) begin
    _zz_io_result_993[1] = _zz_io_result_989[0];
    _zz_io_result_993[0] = (_zz_io_result_989[0] ^ _zz_io_result_989[1]);
  end

  assign _zz_io_result_992 = _zz_io_result_993;
  assign _zz_io_result_994 = ((_zz_io_result_985[0] && _zz_io_result_983[1]) ^ (_zz_io_result_983[0] && _zz_io_result_985[1]));
  always @(*) begin
    _zz_io_result_995[1] = ((_zz_io_result_985[0] && _zz_io_result_983[0]) ^ _zz_io_result_994);
    _zz_io_result_995[0] = ((_zz_io_result_985[1] && _zz_io_result_983[1]) ^ _zz_io_result_994);
  end

  assign _zz_io_result_996 = ((_zz_io_result_986[0] && _zz_io_result_984[1]) ^ (_zz_io_result_984[0] && _zz_io_result_986[1]));
  always @(*) begin
    _zz_io_result_997[1] = ((_zz_io_result_986[0] && _zz_io_result_984[0]) ^ _zz_io_result_996);
    _zz_io_result_997[0] = ((_zz_io_result_986[1] && _zz_io_result_984[1]) ^ _zz_io_result_996);
  end

  always @(*) begin
    _zz_io_result_982[3 : 2] = (_zz_io_result_995 ^ _zz_io_result_992);
    _zz_io_result_982[1 : 0] = (_zz_io_result_997 ^ _zz_io_result_992);
  end

  always @(*) begin
    _zz_io_result_929[7 : 4] = _zz_io_result_982;
    _zz_io_result_929[3 : 0] = _zz_io_result_966;
  end

  assign _zz_io_result_928 = _zz_io_result_929;
  always @(*) begin
    _zz_io_result_999[7] = (_zz_io_result_928[5] ^ _zz_io_result_928[3]);
    _zz_io_result_999[6] = (_zz_io_result_928[7] ^ _zz_io_result_928[3]);
    _zz_io_result_999[5] = (_zz_io_result_928[6] ^ _zz_io_result_928[0]);
    _zz_io_result_999[4] = ((_zz_io_result_928[7] ^ _zz_io_result_928[5]) ^ _zz_io_result_928[3]);
    _zz_io_result_999[3] = ((((_zz_io_result_928[7] ^ _zz_io_result_928[6]) ^ _zz_io_result_928[5]) ^ _zz_io_result_928[4]) ^ _zz_io_result_928[3]);
    _zz_io_result_999[2] = ((((_zz_io_result_928[6] ^ _zz_io_result_928[5]) ^ _zz_io_result_928[3]) ^ _zz_io_result_928[2]) ^ _zz_io_result_928[0]);
    _zz_io_result_999[1] = ((_zz_io_result_928[5] ^ _zz_io_result_928[4]) ^ _zz_io_result_928[1]);
    _zz_io_result_999[0] = ((_zz_io_result_928[6] ^ _zz_io_result_928[4]) ^ _zz_io_result_928[1]);
  end

  assign _zz_io_result_998 = _zz_io_result_999;
  always @(*) begin
    _zz_io_result_925[7] = _zz_io_result_998[7];
    _zz_io_result_925[6] = (! _zz_io_result_998[6]);
    _zz_io_result_925[5] = (! _zz_io_result_998[5]);
    _zz_io_result_925[4] = _zz_io_result_998[4];
    _zz_io_result_925[3] = _zz_io_result_998[3];
    _zz_io_result_925[2] = _zz_io_result_998[2];
    _zz_io_result_925[1] = (! _zz_io_result_998[1]);
    _zz_io_result_925[0] = (! _zz_io_result_998[0]);
  end

  always @(*) begin
    _zz_io_result_923[7 : 0] = _zz_io_result_925;
    _zz_io_result_923[15 : 8] = _zz_io_result_1001;
    _zz_io_result_923[23 : 16] = _zz_io_result_1077;
    _zz_io_result_923[31 : 24] = _zz_io_result_1153;
  end

  assign _zz_io_result_1000 = _zz_io_result_3[15 : 8];
  always @(*) begin
    _zz_io_result_1003[7] = (((((_zz_io_result_1000[7] ^ _zz_io_result_1000[6]) ^ _zz_io_result_1000[5]) ^ _zz_io_result_1000[2]) ^ _zz_io_result_1000[1]) ^ _zz_io_result_1000[0]);
    _zz_io_result_1003[6] = (((_zz_io_result_1000[6] ^ _zz_io_result_1000[5]) ^ _zz_io_result_1000[4]) ^ _zz_io_result_1000[0]);
    _zz_io_result_1003[5] = (((_zz_io_result_1000[6] ^ _zz_io_result_1000[5]) ^ _zz_io_result_1000[1]) ^ _zz_io_result_1000[0]);
    _zz_io_result_1003[4] = (((_zz_io_result_1000[7] ^ _zz_io_result_1000[6]) ^ _zz_io_result_1000[5]) ^ _zz_io_result_1000[0]);
    _zz_io_result_1003[3] = ((((_zz_io_result_1000[7] ^ _zz_io_result_1000[4]) ^ _zz_io_result_1000[3]) ^ _zz_io_result_1000[1]) ^ _zz_io_result_1000[0]);
    _zz_io_result_1003[2] = _zz_io_result_1000[0];
    _zz_io_result_1003[1] = ((_zz_io_result_1000[6] ^ _zz_io_result_1000[5]) ^ _zz_io_result_1000[0]);
    _zz_io_result_1003[0] = ((((_zz_io_result_1000[6] ^ _zz_io_result_1000[3]) ^ _zz_io_result_1000[2]) ^ _zz_io_result_1000[1]) ^ _zz_io_result_1000[0]);
  end

  assign _zz_io_result_1002 = _zz_io_result_1003;
  assign _zz_io_result_1006 = _zz_io_result_1002[7 : 4];
  assign _zz_io_result_1007 = _zz_io_result_1002[3 : 0];
  assign _zz_io_result_1008 = (_zz_io_result_1006 ^ _zz_io_result_1007);
  always @(*) begin
    _zz_io_result_1009[3] = (_zz_io_result_1008[2] ^ _zz_io_result_1008[0]);
    _zz_io_result_1009[2] = (_zz_io_result_1008[3] ^ _zz_io_result_1008[1]);
    _zz_io_result_1009[1] = (_zz_io_result_1008[1] ^ _zz_io_result_1008[0]);
    _zz_io_result_1009[0] = _zz_io_result_1008[0];
  end

  assign _zz_io_result_1011 = _zz_io_result_1006[3 : 2];
  assign _zz_io_result_1012 = _zz_io_result_1006[1 : 0];
  assign _zz_io_result_1013 = _zz_io_result_1007[3 : 2];
  assign _zz_io_result_1014 = _zz_io_result_1007[1 : 0];
  assign _zz_io_result_1015 = (_zz_io_result_1011 ^ _zz_io_result_1012);
  assign _zz_io_result_1016 = (_zz_io_result_1013 ^ _zz_io_result_1014);
  assign _zz_io_result_1018 = ((_zz_io_result_1016[0] && _zz_io_result_1015[1]) ^ (_zz_io_result_1015[0] && _zz_io_result_1016[1]));
  always @(*) begin
    _zz_io_result_1019[1] = ((_zz_io_result_1016[0] && _zz_io_result_1015[0]) ^ _zz_io_result_1018);
    _zz_io_result_1019[0] = ((_zz_io_result_1016[1] && _zz_io_result_1015[1]) ^ _zz_io_result_1018);
  end

  assign _zz_io_result_1017 = _zz_io_result_1019;
  always @(*) begin
    _zz_io_result_1021[1] = _zz_io_result_1017[0];
    _zz_io_result_1021[0] = (_zz_io_result_1017[0] ^ _zz_io_result_1017[1]);
  end

  assign _zz_io_result_1020 = _zz_io_result_1021;
  assign _zz_io_result_1022 = ((_zz_io_result_1013[0] && _zz_io_result_1011[1]) ^ (_zz_io_result_1011[0] && _zz_io_result_1013[1]));
  always @(*) begin
    _zz_io_result_1023[1] = ((_zz_io_result_1013[0] && _zz_io_result_1011[0]) ^ _zz_io_result_1022);
    _zz_io_result_1023[0] = ((_zz_io_result_1013[1] && _zz_io_result_1011[1]) ^ _zz_io_result_1022);
  end

  assign _zz_io_result_1024 = ((_zz_io_result_1014[0] && _zz_io_result_1012[1]) ^ (_zz_io_result_1012[0] && _zz_io_result_1014[1]));
  always @(*) begin
    _zz_io_result_1025[1] = ((_zz_io_result_1014[0] && _zz_io_result_1012[0]) ^ _zz_io_result_1024);
    _zz_io_result_1025[0] = ((_zz_io_result_1014[1] && _zz_io_result_1012[1]) ^ _zz_io_result_1024);
  end

  always @(*) begin
    _zz_io_result_1010[3 : 2] = (_zz_io_result_1023 ^ _zz_io_result_1020);
    _zz_io_result_1010[1 : 0] = (_zz_io_result_1025 ^ _zz_io_result_1020);
  end

  assign _zz_io_result_1026 = (_zz_io_result_1009 ^ _zz_io_result_1010);
  assign _zz_io_result_1029 = _zz_io_result_1026[3 : 2];
  assign _zz_io_result_1030 = _zz_io_result_1026[1 : 0];
  assign _zz_io_result_1031 = (_zz_io_result_1029 ^ _zz_io_result_1030);
  always @(*) begin
    _zz_io_result_1032[1] = _zz_io_result_1031[1];
    _zz_io_result_1032[0] = (_zz_io_result_1031[0] ^ _zz_io_result_1031[1]);
  end

  assign _zz_io_result_1033 = ((_zz_io_result_1030[0] && _zz_io_result_1029[1]) ^ (_zz_io_result_1029[0] && _zz_io_result_1030[1]));
  always @(*) begin
    _zz_io_result_1034[1] = ((_zz_io_result_1030[0] && _zz_io_result_1029[0]) ^ _zz_io_result_1033);
    _zz_io_result_1034[0] = ((_zz_io_result_1030[1] && _zz_io_result_1029[1]) ^ _zz_io_result_1033);
  end

  assign _zz_io_result_1035 = (_zz_io_result_1032 ^ _zz_io_result_1034);
  always @(*) begin
    _zz_io_result_1037[1] = _zz_io_result_1035[0];
    _zz_io_result_1037[0] = _zz_io_result_1035[1];
  end

  assign _zz_io_result_1036 = _zz_io_result_1037;
  assign _zz_io_result_1038 = ((_zz_io_result_1036[0] && _zz_io_result_1029[1]) ^ (_zz_io_result_1029[0] && _zz_io_result_1036[1]));
  always @(*) begin
    _zz_io_result_1039[1] = ((_zz_io_result_1036[0] && _zz_io_result_1029[0]) ^ _zz_io_result_1038);
    _zz_io_result_1039[0] = ((_zz_io_result_1036[1] && _zz_io_result_1029[1]) ^ _zz_io_result_1038);
  end

  assign _zz_io_result_1040 = ((_zz_io_result_1036[0] && _zz_io_result_1030[1]) ^ (_zz_io_result_1030[0] && _zz_io_result_1036[1]));
  always @(*) begin
    _zz_io_result_1041[1] = ((_zz_io_result_1036[0] && _zz_io_result_1030[0]) ^ _zz_io_result_1040);
    _zz_io_result_1041[0] = ((_zz_io_result_1036[1] && _zz_io_result_1030[1]) ^ _zz_io_result_1040);
  end

  always @(*) begin
    _zz_io_result_1028[3 : 2] = _zz_io_result_1041;
    _zz_io_result_1028[1 : 0] = _zz_io_result_1039;
  end

  assign _zz_io_result_1027 = _zz_io_result_1028;
  assign _zz_io_result_1043 = _zz_io_result_1006[3 : 2];
  assign _zz_io_result_1044 = _zz_io_result_1006[1 : 0];
  assign _zz_io_result_1045 = _zz_io_result_1027[3 : 2];
  assign _zz_io_result_1046 = _zz_io_result_1027[1 : 0];
  assign _zz_io_result_1047 = (_zz_io_result_1043 ^ _zz_io_result_1044);
  assign _zz_io_result_1048 = (_zz_io_result_1045 ^ _zz_io_result_1046);
  assign _zz_io_result_1050 = ((_zz_io_result_1048[0] && _zz_io_result_1047[1]) ^ (_zz_io_result_1047[0] && _zz_io_result_1048[1]));
  always @(*) begin
    _zz_io_result_1051[1] = ((_zz_io_result_1048[0] && _zz_io_result_1047[0]) ^ _zz_io_result_1050);
    _zz_io_result_1051[0] = ((_zz_io_result_1048[1] && _zz_io_result_1047[1]) ^ _zz_io_result_1050);
  end

  assign _zz_io_result_1049 = _zz_io_result_1051;
  always @(*) begin
    _zz_io_result_1053[1] = _zz_io_result_1049[0];
    _zz_io_result_1053[0] = (_zz_io_result_1049[0] ^ _zz_io_result_1049[1]);
  end

  assign _zz_io_result_1052 = _zz_io_result_1053;
  assign _zz_io_result_1054 = ((_zz_io_result_1045[0] && _zz_io_result_1043[1]) ^ (_zz_io_result_1043[0] && _zz_io_result_1045[1]));
  always @(*) begin
    _zz_io_result_1055[1] = ((_zz_io_result_1045[0] && _zz_io_result_1043[0]) ^ _zz_io_result_1054);
    _zz_io_result_1055[0] = ((_zz_io_result_1045[1] && _zz_io_result_1043[1]) ^ _zz_io_result_1054);
  end

  assign _zz_io_result_1056 = ((_zz_io_result_1046[0] && _zz_io_result_1044[1]) ^ (_zz_io_result_1044[0] && _zz_io_result_1046[1]));
  always @(*) begin
    _zz_io_result_1057[1] = ((_zz_io_result_1046[0] && _zz_io_result_1044[0]) ^ _zz_io_result_1056);
    _zz_io_result_1057[0] = ((_zz_io_result_1046[1] && _zz_io_result_1044[1]) ^ _zz_io_result_1056);
  end

  always @(*) begin
    _zz_io_result_1042[3 : 2] = (_zz_io_result_1055 ^ _zz_io_result_1052);
    _zz_io_result_1042[1 : 0] = (_zz_io_result_1057 ^ _zz_io_result_1052);
  end

  assign _zz_io_result_1059 = _zz_io_result_1007[3 : 2];
  assign _zz_io_result_1060 = _zz_io_result_1007[1 : 0];
  assign _zz_io_result_1061 = _zz_io_result_1027[3 : 2];
  assign _zz_io_result_1062 = _zz_io_result_1027[1 : 0];
  assign _zz_io_result_1063 = (_zz_io_result_1059 ^ _zz_io_result_1060);
  assign _zz_io_result_1064 = (_zz_io_result_1061 ^ _zz_io_result_1062);
  assign _zz_io_result_1066 = ((_zz_io_result_1064[0] && _zz_io_result_1063[1]) ^ (_zz_io_result_1063[0] && _zz_io_result_1064[1]));
  always @(*) begin
    _zz_io_result_1067[1] = ((_zz_io_result_1064[0] && _zz_io_result_1063[0]) ^ _zz_io_result_1066);
    _zz_io_result_1067[0] = ((_zz_io_result_1064[1] && _zz_io_result_1063[1]) ^ _zz_io_result_1066);
  end

  assign _zz_io_result_1065 = _zz_io_result_1067;
  always @(*) begin
    _zz_io_result_1069[1] = _zz_io_result_1065[0];
    _zz_io_result_1069[0] = (_zz_io_result_1065[0] ^ _zz_io_result_1065[1]);
  end

  assign _zz_io_result_1068 = _zz_io_result_1069;
  assign _zz_io_result_1070 = ((_zz_io_result_1061[0] && _zz_io_result_1059[1]) ^ (_zz_io_result_1059[0] && _zz_io_result_1061[1]));
  always @(*) begin
    _zz_io_result_1071[1] = ((_zz_io_result_1061[0] && _zz_io_result_1059[0]) ^ _zz_io_result_1070);
    _zz_io_result_1071[0] = ((_zz_io_result_1061[1] && _zz_io_result_1059[1]) ^ _zz_io_result_1070);
  end

  assign _zz_io_result_1072 = ((_zz_io_result_1062[0] && _zz_io_result_1060[1]) ^ (_zz_io_result_1060[0] && _zz_io_result_1062[1]));
  always @(*) begin
    _zz_io_result_1073[1] = ((_zz_io_result_1062[0] && _zz_io_result_1060[0]) ^ _zz_io_result_1072);
    _zz_io_result_1073[0] = ((_zz_io_result_1062[1] && _zz_io_result_1060[1]) ^ _zz_io_result_1072);
  end

  always @(*) begin
    _zz_io_result_1058[3 : 2] = (_zz_io_result_1071 ^ _zz_io_result_1068);
    _zz_io_result_1058[1 : 0] = (_zz_io_result_1073 ^ _zz_io_result_1068);
  end

  always @(*) begin
    _zz_io_result_1005[7 : 4] = _zz_io_result_1058;
    _zz_io_result_1005[3 : 0] = _zz_io_result_1042;
  end

  assign _zz_io_result_1004 = _zz_io_result_1005;
  always @(*) begin
    _zz_io_result_1075[7] = (_zz_io_result_1004[5] ^ _zz_io_result_1004[3]);
    _zz_io_result_1075[6] = (_zz_io_result_1004[7] ^ _zz_io_result_1004[3]);
    _zz_io_result_1075[5] = (_zz_io_result_1004[6] ^ _zz_io_result_1004[0]);
    _zz_io_result_1075[4] = ((_zz_io_result_1004[7] ^ _zz_io_result_1004[5]) ^ _zz_io_result_1004[3]);
    _zz_io_result_1075[3] = ((((_zz_io_result_1004[7] ^ _zz_io_result_1004[6]) ^ _zz_io_result_1004[5]) ^ _zz_io_result_1004[4]) ^ _zz_io_result_1004[3]);
    _zz_io_result_1075[2] = ((((_zz_io_result_1004[6] ^ _zz_io_result_1004[5]) ^ _zz_io_result_1004[3]) ^ _zz_io_result_1004[2]) ^ _zz_io_result_1004[0]);
    _zz_io_result_1075[1] = ((_zz_io_result_1004[5] ^ _zz_io_result_1004[4]) ^ _zz_io_result_1004[1]);
    _zz_io_result_1075[0] = ((_zz_io_result_1004[6] ^ _zz_io_result_1004[4]) ^ _zz_io_result_1004[1]);
  end

  assign _zz_io_result_1074 = _zz_io_result_1075;
  always @(*) begin
    _zz_io_result_1001[7] = _zz_io_result_1074[7];
    _zz_io_result_1001[6] = (! _zz_io_result_1074[6]);
    _zz_io_result_1001[5] = (! _zz_io_result_1074[5]);
    _zz_io_result_1001[4] = _zz_io_result_1074[4];
    _zz_io_result_1001[3] = _zz_io_result_1074[3];
    _zz_io_result_1001[2] = _zz_io_result_1074[2];
    _zz_io_result_1001[1] = (! _zz_io_result_1074[1]);
    _zz_io_result_1001[0] = (! _zz_io_result_1074[0]);
  end

  assign _zz_io_result_1076 = _zz_io_result_3[23 : 16];
  always @(*) begin
    _zz_io_result_1079[7] = (((((_zz_io_result_1076[7] ^ _zz_io_result_1076[6]) ^ _zz_io_result_1076[5]) ^ _zz_io_result_1076[2]) ^ _zz_io_result_1076[1]) ^ _zz_io_result_1076[0]);
    _zz_io_result_1079[6] = (((_zz_io_result_1076[6] ^ _zz_io_result_1076[5]) ^ _zz_io_result_1076[4]) ^ _zz_io_result_1076[0]);
    _zz_io_result_1079[5] = (((_zz_io_result_1076[6] ^ _zz_io_result_1076[5]) ^ _zz_io_result_1076[1]) ^ _zz_io_result_1076[0]);
    _zz_io_result_1079[4] = (((_zz_io_result_1076[7] ^ _zz_io_result_1076[6]) ^ _zz_io_result_1076[5]) ^ _zz_io_result_1076[0]);
    _zz_io_result_1079[3] = ((((_zz_io_result_1076[7] ^ _zz_io_result_1076[4]) ^ _zz_io_result_1076[3]) ^ _zz_io_result_1076[1]) ^ _zz_io_result_1076[0]);
    _zz_io_result_1079[2] = _zz_io_result_1076[0];
    _zz_io_result_1079[1] = ((_zz_io_result_1076[6] ^ _zz_io_result_1076[5]) ^ _zz_io_result_1076[0]);
    _zz_io_result_1079[0] = ((((_zz_io_result_1076[6] ^ _zz_io_result_1076[3]) ^ _zz_io_result_1076[2]) ^ _zz_io_result_1076[1]) ^ _zz_io_result_1076[0]);
  end

  assign _zz_io_result_1078 = _zz_io_result_1079;
  assign _zz_io_result_1082 = _zz_io_result_1078[7 : 4];
  assign _zz_io_result_1083 = _zz_io_result_1078[3 : 0];
  assign _zz_io_result_1084 = (_zz_io_result_1082 ^ _zz_io_result_1083);
  always @(*) begin
    _zz_io_result_1085[3] = (_zz_io_result_1084[2] ^ _zz_io_result_1084[0]);
    _zz_io_result_1085[2] = (_zz_io_result_1084[3] ^ _zz_io_result_1084[1]);
    _zz_io_result_1085[1] = (_zz_io_result_1084[1] ^ _zz_io_result_1084[0]);
    _zz_io_result_1085[0] = _zz_io_result_1084[0];
  end

  assign _zz_io_result_1087 = _zz_io_result_1082[3 : 2];
  assign _zz_io_result_1088 = _zz_io_result_1082[1 : 0];
  assign _zz_io_result_1089 = _zz_io_result_1083[3 : 2];
  assign _zz_io_result_1090 = _zz_io_result_1083[1 : 0];
  assign _zz_io_result_1091 = (_zz_io_result_1087 ^ _zz_io_result_1088);
  assign _zz_io_result_1092 = (_zz_io_result_1089 ^ _zz_io_result_1090);
  assign _zz_io_result_1094 = ((_zz_io_result_1092[0] && _zz_io_result_1091[1]) ^ (_zz_io_result_1091[0] && _zz_io_result_1092[1]));
  always @(*) begin
    _zz_io_result_1095[1] = ((_zz_io_result_1092[0] && _zz_io_result_1091[0]) ^ _zz_io_result_1094);
    _zz_io_result_1095[0] = ((_zz_io_result_1092[1] && _zz_io_result_1091[1]) ^ _zz_io_result_1094);
  end

  assign _zz_io_result_1093 = _zz_io_result_1095;
  always @(*) begin
    _zz_io_result_1097[1] = _zz_io_result_1093[0];
    _zz_io_result_1097[0] = (_zz_io_result_1093[0] ^ _zz_io_result_1093[1]);
  end

  assign _zz_io_result_1096 = _zz_io_result_1097;
  assign _zz_io_result_1098 = ((_zz_io_result_1089[0] && _zz_io_result_1087[1]) ^ (_zz_io_result_1087[0] && _zz_io_result_1089[1]));
  always @(*) begin
    _zz_io_result_1099[1] = ((_zz_io_result_1089[0] && _zz_io_result_1087[0]) ^ _zz_io_result_1098);
    _zz_io_result_1099[0] = ((_zz_io_result_1089[1] && _zz_io_result_1087[1]) ^ _zz_io_result_1098);
  end

  assign _zz_io_result_1100 = ((_zz_io_result_1090[0] && _zz_io_result_1088[1]) ^ (_zz_io_result_1088[0] && _zz_io_result_1090[1]));
  always @(*) begin
    _zz_io_result_1101[1] = ((_zz_io_result_1090[0] && _zz_io_result_1088[0]) ^ _zz_io_result_1100);
    _zz_io_result_1101[0] = ((_zz_io_result_1090[1] && _zz_io_result_1088[1]) ^ _zz_io_result_1100);
  end

  always @(*) begin
    _zz_io_result_1086[3 : 2] = (_zz_io_result_1099 ^ _zz_io_result_1096);
    _zz_io_result_1086[1 : 0] = (_zz_io_result_1101 ^ _zz_io_result_1096);
  end

  assign _zz_io_result_1102 = (_zz_io_result_1085 ^ _zz_io_result_1086);
  assign _zz_io_result_1105 = _zz_io_result_1102[3 : 2];
  assign _zz_io_result_1106 = _zz_io_result_1102[1 : 0];
  assign _zz_io_result_1107 = (_zz_io_result_1105 ^ _zz_io_result_1106);
  always @(*) begin
    _zz_io_result_1108[1] = _zz_io_result_1107[1];
    _zz_io_result_1108[0] = (_zz_io_result_1107[0] ^ _zz_io_result_1107[1]);
  end

  assign _zz_io_result_1109 = ((_zz_io_result_1106[0] && _zz_io_result_1105[1]) ^ (_zz_io_result_1105[0] && _zz_io_result_1106[1]));
  always @(*) begin
    _zz_io_result_1110[1] = ((_zz_io_result_1106[0] && _zz_io_result_1105[0]) ^ _zz_io_result_1109);
    _zz_io_result_1110[0] = ((_zz_io_result_1106[1] && _zz_io_result_1105[1]) ^ _zz_io_result_1109);
  end

  assign _zz_io_result_1111 = (_zz_io_result_1108 ^ _zz_io_result_1110);
  always @(*) begin
    _zz_io_result_1113[1] = _zz_io_result_1111[0];
    _zz_io_result_1113[0] = _zz_io_result_1111[1];
  end

  assign _zz_io_result_1112 = _zz_io_result_1113;
  assign _zz_io_result_1114 = ((_zz_io_result_1112[0] && _zz_io_result_1105[1]) ^ (_zz_io_result_1105[0] && _zz_io_result_1112[1]));
  always @(*) begin
    _zz_io_result_1115[1] = ((_zz_io_result_1112[0] && _zz_io_result_1105[0]) ^ _zz_io_result_1114);
    _zz_io_result_1115[0] = ((_zz_io_result_1112[1] && _zz_io_result_1105[1]) ^ _zz_io_result_1114);
  end

  assign _zz_io_result_1116 = ((_zz_io_result_1112[0] && _zz_io_result_1106[1]) ^ (_zz_io_result_1106[0] && _zz_io_result_1112[1]));
  always @(*) begin
    _zz_io_result_1117[1] = ((_zz_io_result_1112[0] && _zz_io_result_1106[0]) ^ _zz_io_result_1116);
    _zz_io_result_1117[0] = ((_zz_io_result_1112[1] && _zz_io_result_1106[1]) ^ _zz_io_result_1116);
  end

  always @(*) begin
    _zz_io_result_1104[3 : 2] = _zz_io_result_1117;
    _zz_io_result_1104[1 : 0] = _zz_io_result_1115;
  end

  assign _zz_io_result_1103 = _zz_io_result_1104;
  assign _zz_io_result_1119 = _zz_io_result_1082[3 : 2];
  assign _zz_io_result_1120 = _zz_io_result_1082[1 : 0];
  assign _zz_io_result_1121 = _zz_io_result_1103[3 : 2];
  assign _zz_io_result_1122 = _zz_io_result_1103[1 : 0];
  assign _zz_io_result_1123 = (_zz_io_result_1119 ^ _zz_io_result_1120);
  assign _zz_io_result_1124 = (_zz_io_result_1121 ^ _zz_io_result_1122);
  assign _zz_io_result_1126 = ((_zz_io_result_1124[0] && _zz_io_result_1123[1]) ^ (_zz_io_result_1123[0] && _zz_io_result_1124[1]));
  always @(*) begin
    _zz_io_result_1127[1] = ((_zz_io_result_1124[0] && _zz_io_result_1123[0]) ^ _zz_io_result_1126);
    _zz_io_result_1127[0] = ((_zz_io_result_1124[1] && _zz_io_result_1123[1]) ^ _zz_io_result_1126);
  end

  assign _zz_io_result_1125 = _zz_io_result_1127;
  always @(*) begin
    _zz_io_result_1129[1] = _zz_io_result_1125[0];
    _zz_io_result_1129[0] = (_zz_io_result_1125[0] ^ _zz_io_result_1125[1]);
  end

  assign _zz_io_result_1128 = _zz_io_result_1129;
  assign _zz_io_result_1130 = ((_zz_io_result_1121[0] && _zz_io_result_1119[1]) ^ (_zz_io_result_1119[0] && _zz_io_result_1121[1]));
  always @(*) begin
    _zz_io_result_1131[1] = ((_zz_io_result_1121[0] && _zz_io_result_1119[0]) ^ _zz_io_result_1130);
    _zz_io_result_1131[0] = ((_zz_io_result_1121[1] && _zz_io_result_1119[1]) ^ _zz_io_result_1130);
  end

  assign _zz_io_result_1132 = ((_zz_io_result_1122[0] && _zz_io_result_1120[1]) ^ (_zz_io_result_1120[0] && _zz_io_result_1122[1]));
  always @(*) begin
    _zz_io_result_1133[1] = ((_zz_io_result_1122[0] && _zz_io_result_1120[0]) ^ _zz_io_result_1132);
    _zz_io_result_1133[0] = ((_zz_io_result_1122[1] && _zz_io_result_1120[1]) ^ _zz_io_result_1132);
  end

  always @(*) begin
    _zz_io_result_1118[3 : 2] = (_zz_io_result_1131 ^ _zz_io_result_1128);
    _zz_io_result_1118[1 : 0] = (_zz_io_result_1133 ^ _zz_io_result_1128);
  end

  assign _zz_io_result_1135 = _zz_io_result_1083[3 : 2];
  assign _zz_io_result_1136 = _zz_io_result_1083[1 : 0];
  assign _zz_io_result_1137 = _zz_io_result_1103[3 : 2];
  assign _zz_io_result_1138 = _zz_io_result_1103[1 : 0];
  assign _zz_io_result_1139 = (_zz_io_result_1135 ^ _zz_io_result_1136);
  assign _zz_io_result_1140 = (_zz_io_result_1137 ^ _zz_io_result_1138);
  assign _zz_io_result_1142 = ((_zz_io_result_1140[0] && _zz_io_result_1139[1]) ^ (_zz_io_result_1139[0] && _zz_io_result_1140[1]));
  always @(*) begin
    _zz_io_result_1143[1] = ((_zz_io_result_1140[0] && _zz_io_result_1139[0]) ^ _zz_io_result_1142);
    _zz_io_result_1143[0] = ((_zz_io_result_1140[1] && _zz_io_result_1139[1]) ^ _zz_io_result_1142);
  end

  assign _zz_io_result_1141 = _zz_io_result_1143;
  always @(*) begin
    _zz_io_result_1145[1] = _zz_io_result_1141[0];
    _zz_io_result_1145[0] = (_zz_io_result_1141[0] ^ _zz_io_result_1141[1]);
  end

  assign _zz_io_result_1144 = _zz_io_result_1145;
  assign _zz_io_result_1146 = ((_zz_io_result_1137[0] && _zz_io_result_1135[1]) ^ (_zz_io_result_1135[0] && _zz_io_result_1137[1]));
  always @(*) begin
    _zz_io_result_1147[1] = ((_zz_io_result_1137[0] && _zz_io_result_1135[0]) ^ _zz_io_result_1146);
    _zz_io_result_1147[0] = ((_zz_io_result_1137[1] && _zz_io_result_1135[1]) ^ _zz_io_result_1146);
  end

  assign _zz_io_result_1148 = ((_zz_io_result_1138[0] && _zz_io_result_1136[1]) ^ (_zz_io_result_1136[0] && _zz_io_result_1138[1]));
  always @(*) begin
    _zz_io_result_1149[1] = ((_zz_io_result_1138[0] && _zz_io_result_1136[0]) ^ _zz_io_result_1148);
    _zz_io_result_1149[0] = ((_zz_io_result_1138[1] && _zz_io_result_1136[1]) ^ _zz_io_result_1148);
  end

  always @(*) begin
    _zz_io_result_1134[3 : 2] = (_zz_io_result_1147 ^ _zz_io_result_1144);
    _zz_io_result_1134[1 : 0] = (_zz_io_result_1149 ^ _zz_io_result_1144);
  end

  always @(*) begin
    _zz_io_result_1081[7 : 4] = _zz_io_result_1134;
    _zz_io_result_1081[3 : 0] = _zz_io_result_1118;
  end

  assign _zz_io_result_1080 = _zz_io_result_1081;
  always @(*) begin
    _zz_io_result_1151[7] = (_zz_io_result_1080[5] ^ _zz_io_result_1080[3]);
    _zz_io_result_1151[6] = (_zz_io_result_1080[7] ^ _zz_io_result_1080[3]);
    _zz_io_result_1151[5] = (_zz_io_result_1080[6] ^ _zz_io_result_1080[0]);
    _zz_io_result_1151[4] = ((_zz_io_result_1080[7] ^ _zz_io_result_1080[5]) ^ _zz_io_result_1080[3]);
    _zz_io_result_1151[3] = ((((_zz_io_result_1080[7] ^ _zz_io_result_1080[6]) ^ _zz_io_result_1080[5]) ^ _zz_io_result_1080[4]) ^ _zz_io_result_1080[3]);
    _zz_io_result_1151[2] = ((((_zz_io_result_1080[6] ^ _zz_io_result_1080[5]) ^ _zz_io_result_1080[3]) ^ _zz_io_result_1080[2]) ^ _zz_io_result_1080[0]);
    _zz_io_result_1151[1] = ((_zz_io_result_1080[5] ^ _zz_io_result_1080[4]) ^ _zz_io_result_1080[1]);
    _zz_io_result_1151[0] = ((_zz_io_result_1080[6] ^ _zz_io_result_1080[4]) ^ _zz_io_result_1080[1]);
  end

  assign _zz_io_result_1150 = _zz_io_result_1151;
  always @(*) begin
    _zz_io_result_1077[7] = _zz_io_result_1150[7];
    _zz_io_result_1077[6] = (! _zz_io_result_1150[6]);
    _zz_io_result_1077[5] = (! _zz_io_result_1150[5]);
    _zz_io_result_1077[4] = _zz_io_result_1150[4];
    _zz_io_result_1077[3] = _zz_io_result_1150[3];
    _zz_io_result_1077[2] = _zz_io_result_1150[2];
    _zz_io_result_1077[1] = (! _zz_io_result_1150[1]);
    _zz_io_result_1077[0] = (! _zz_io_result_1150[0]);
  end

  assign _zz_io_result_1152 = _zz_io_result_3[31 : 24];
  always @(*) begin
    _zz_io_result_1155[7] = (((((_zz_io_result_1152[7] ^ _zz_io_result_1152[6]) ^ _zz_io_result_1152[5]) ^ _zz_io_result_1152[2]) ^ _zz_io_result_1152[1]) ^ _zz_io_result_1152[0]);
    _zz_io_result_1155[6] = (((_zz_io_result_1152[6] ^ _zz_io_result_1152[5]) ^ _zz_io_result_1152[4]) ^ _zz_io_result_1152[0]);
    _zz_io_result_1155[5] = (((_zz_io_result_1152[6] ^ _zz_io_result_1152[5]) ^ _zz_io_result_1152[1]) ^ _zz_io_result_1152[0]);
    _zz_io_result_1155[4] = (((_zz_io_result_1152[7] ^ _zz_io_result_1152[6]) ^ _zz_io_result_1152[5]) ^ _zz_io_result_1152[0]);
    _zz_io_result_1155[3] = ((((_zz_io_result_1152[7] ^ _zz_io_result_1152[4]) ^ _zz_io_result_1152[3]) ^ _zz_io_result_1152[1]) ^ _zz_io_result_1152[0]);
    _zz_io_result_1155[2] = _zz_io_result_1152[0];
    _zz_io_result_1155[1] = ((_zz_io_result_1152[6] ^ _zz_io_result_1152[5]) ^ _zz_io_result_1152[0]);
    _zz_io_result_1155[0] = ((((_zz_io_result_1152[6] ^ _zz_io_result_1152[3]) ^ _zz_io_result_1152[2]) ^ _zz_io_result_1152[1]) ^ _zz_io_result_1152[0]);
  end

  assign _zz_io_result_1154 = _zz_io_result_1155;
  assign _zz_io_result_1158 = _zz_io_result_1154[7 : 4];
  assign _zz_io_result_1159 = _zz_io_result_1154[3 : 0];
  assign _zz_io_result_1160 = (_zz_io_result_1158 ^ _zz_io_result_1159);
  always @(*) begin
    _zz_io_result_1161[3] = (_zz_io_result_1160[2] ^ _zz_io_result_1160[0]);
    _zz_io_result_1161[2] = (_zz_io_result_1160[3] ^ _zz_io_result_1160[1]);
    _zz_io_result_1161[1] = (_zz_io_result_1160[1] ^ _zz_io_result_1160[0]);
    _zz_io_result_1161[0] = _zz_io_result_1160[0];
  end

  assign _zz_io_result_1163 = _zz_io_result_1158[3 : 2];
  assign _zz_io_result_1164 = _zz_io_result_1158[1 : 0];
  assign _zz_io_result_1165 = _zz_io_result_1159[3 : 2];
  assign _zz_io_result_1166 = _zz_io_result_1159[1 : 0];
  assign _zz_io_result_1167 = (_zz_io_result_1163 ^ _zz_io_result_1164);
  assign _zz_io_result_1168 = (_zz_io_result_1165 ^ _zz_io_result_1166);
  assign _zz_io_result_1170 = ((_zz_io_result_1168[0] && _zz_io_result_1167[1]) ^ (_zz_io_result_1167[0] && _zz_io_result_1168[1]));
  always @(*) begin
    _zz_io_result_1171[1] = ((_zz_io_result_1168[0] && _zz_io_result_1167[0]) ^ _zz_io_result_1170);
    _zz_io_result_1171[0] = ((_zz_io_result_1168[1] && _zz_io_result_1167[1]) ^ _zz_io_result_1170);
  end

  assign _zz_io_result_1169 = _zz_io_result_1171;
  always @(*) begin
    _zz_io_result_1173[1] = _zz_io_result_1169[0];
    _zz_io_result_1173[0] = (_zz_io_result_1169[0] ^ _zz_io_result_1169[1]);
  end

  assign _zz_io_result_1172 = _zz_io_result_1173;
  assign _zz_io_result_1174 = ((_zz_io_result_1165[0] && _zz_io_result_1163[1]) ^ (_zz_io_result_1163[0] && _zz_io_result_1165[1]));
  always @(*) begin
    _zz_io_result_1175[1] = ((_zz_io_result_1165[0] && _zz_io_result_1163[0]) ^ _zz_io_result_1174);
    _zz_io_result_1175[0] = ((_zz_io_result_1165[1] && _zz_io_result_1163[1]) ^ _zz_io_result_1174);
  end

  assign _zz_io_result_1176 = ((_zz_io_result_1166[0] && _zz_io_result_1164[1]) ^ (_zz_io_result_1164[0] && _zz_io_result_1166[1]));
  always @(*) begin
    _zz_io_result_1177[1] = ((_zz_io_result_1166[0] && _zz_io_result_1164[0]) ^ _zz_io_result_1176);
    _zz_io_result_1177[0] = ((_zz_io_result_1166[1] && _zz_io_result_1164[1]) ^ _zz_io_result_1176);
  end

  always @(*) begin
    _zz_io_result_1162[3 : 2] = (_zz_io_result_1175 ^ _zz_io_result_1172);
    _zz_io_result_1162[1 : 0] = (_zz_io_result_1177 ^ _zz_io_result_1172);
  end

  assign _zz_io_result_1178 = (_zz_io_result_1161 ^ _zz_io_result_1162);
  assign _zz_io_result_1181 = _zz_io_result_1178[3 : 2];
  assign _zz_io_result_1182 = _zz_io_result_1178[1 : 0];
  assign _zz_io_result_1183 = (_zz_io_result_1181 ^ _zz_io_result_1182);
  always @(*) begin
    _zz_io_result_1184[1] = _zz_io_result_1183[1];
    _zz_io_result_1184[0] = (_zz_io_result_1183[0] ^ _zz_io_result_1183[1]);
  end

  assign _zz_io_result_1185 = ((_zz_io_result_1182[0] && _zz_io_result_1181[1]) ^ (_zz_io_result_1181[0] && _zz_io_result_1182[1]));
  always @(*) begin
    _zz_io_result_1186[1] = ((_zz_io_result_1182[0] && _zz_io_result_1181[0]) ^ _zz_io_result_1185);
    _zz_io_result_1186[0] = ((_zz_io_result_1182[1] && _zz_io_result_1181[1]) ^ _zz_io_result_1185);
  end

  assign _zz_io_result_1187 = (_zz_io_result_1184 ^ _zz_io_result_1186);
  always @(*) begin
    _zz_io_result_1189[1] = _zz_io_result_1187[0];
    _zz_io_result_1189[0] = _zz_io_result_1187[1];
  end

  assign _zz_io_result_1188 = _zz_io_result_1189;
  assign _zz_io_result_1190 = ((_zz_io_result_1188[0] && _zz_io_result_1181[1]) ^ (_zz_io_result_1181[0] && _zz_io_result_1188[1]));
  always @(*) begin
    _zz_io_result_1191[1] = ((_zz_io_result_1188[0] && _zz_io_result_1181[0]) ^ _zz_io_result_1190);
    _zz_io_result_1191[0] = ((_zz_io_result_1188[1] && _zz_io_result_1181[1]) ^ _zz_io_result_1190);
  end

  assign _zz_io_result_1192 = ((_zz_io_result_1188[0] && _zz_io_result_1182[1]) ^ (_zz_io_result_1182[0] && _zz_io_result_1188[1]));
  always @(*) begin
    _zz_io_result_1193[1] = ((_zz_io_result_1188[0] && _zz_io_result_1182[0]) ^ _zz_io_result_1192);
    _zz_io_result_1193[0] = ((_zz_io_result_1188[1] && _zz_io_result_1182[1]) ^ _zz_io_result_1192);
  end

  always @(*) begin
    _zz_io_result_1180[3 : 2] = _zz_io_result_1193;
    _zz_io_result_1180[1 : 0] = _zz_io_result_1191;
  end

  assign _zz_io_result_1179 = _zz_io_result_1180;
  assign _zz_io_result_1195 = _zz_io_result_1158[3 : 2];
  assign _zz_io_result_1196 = _zz_io_result_1158[1 : 0];
  assign _zz_io_result_1197 = _zz_io_result_1179[3 : 2];
  assign _zz_io_result_1198 = _zz_io_result_1179[1 : 0];
  assign _zz_io_result_1199 = (_zz_io_result_1195 ^ _zz_io_result_1196);
  assign _zz_io_result_1200 = (_zz_io_result_1197 ^ _zz_io_result_1198);
  assign _zz_io_result_1202 = ((_zz_io_result_1200[0] && _zz_io_result_1199[1]) ^ (_zz_io_result_1199[0] && _zz_io_result_1200[1]));
  always @(*) begin
    _zz_io_result_1203[1] = ((_zz_io_result_1200[0] && _zz_io_result_1199[0]) ^ _zz_io_result_1202);
    _zz_io_result_1203[0] = ((_zz_io_result_1200[1] && _zz_io_result_1199[1]) ^ _zz_io_result_1202);
  end

  assign _zz_io_result_1201 = _zz_io_result_1203;
  always @(*) begin
    _zz_io_result_1205[1] = _zz_io_result_1201[0];
    _zz_io_result_1205[0] = (_zz_io_result_1201[0] ^ _zz_io_result_1201[1]);
  end

  assign _zz_io_result_1204 = _zz_io_result_1205;
  assign _zz_io_result_1206 = ((_zz_io_result_1197[0] && _zz_io_result_1195[1]) ^ (_zz_io_result_1195[0] && _zz_io_result_1197[1]));
  always @(*) begin
    _zz_io_result_1207[1] = ((_zz_io_result_1197[0] && _zz_io_result_1195[0]) ^ _zz_io_result_1206);
    _zz_io_result_1207[0] = ((_zz_io_result_1197[1] && _zz_io_result_1195[1]) ^ _zz_io_result_1206);
  end

  assign _zz_io_result_1208 = ((_zz_io_result_1198[0] && _zz_io_result_1196[1]) ^ (_zz_io_result_1196[0] && _zz_io_result_1198[1]));
  always @(*) begin
    _zz_io_result_1209[1] = ((_zz_io_result_1198[0] && _zz_io_result_1196[0]) ^ _zz_io_result_1208);
    _zz_io_result_1209[0] = ((_zz_io_result_1198[1] && _zz_io_result_1196[1]) ^ _zz_io_result_1208);
  end

  always @(*) begin
    _zz_io_result_1194[3 : 2] = (_zz_io_result_1207 ^ _zz_io_result_1204);
    _zz_io_result_1194[1 : 0] = (_zz_io_result_1209 ^ _zz_io_result_1204);
  end

  assign _zz_io_result_1211 = _zz_io_result_1159[3 : 2];
  assign _zz_io_result_1212 = _zz_io_result_1159[1 : 0];
  assign _zz_io_result_1213 = _zz_io_result_1179[3 : 2];
  assign _zz_io_result_1214 = _zz_io_result_1179[1 : 0];
  assign _zz_io_result_1215 = (_zz_io_result_1211 ^ _zz_io_result_1212);
  assign _zz_io_result_1216 = (_zz_io_result_1213 ^ _zz_io_result_1214);
  assign _zz_io_result_1218 = ((_zz_io_result_1216[0] && _zz_io_result_1215[1]) ^ (_zz_io_result_1215[0] && _zz_io_result_1216[1]));
  always @(*) begin
    _zz_io_result_1219[1] = ((_zz_io_result_1216[0] && _zz_io_result_1215[0]) ^ _zz_io_result_1218);
    _zz_io_result_1219[0] = ((_zz_io_result_1216[1] && _zz_io_result_1215[1]) ^ _zz_io_result_1218);
  end

  assign _zz_io_result_1217 = _zz_io_result_1219;
  always @(*) begin
    _zz_io_result_1221[1] = _zz_io_result_1217[0];
    _zz_io_result_1221[0] = (_zz_io_result_1217[0] ^ _zz_io_result_1217[1]);
  end

  assign _zz_io_result_1220 = _zz_io_result_1221;
  assign _zz_io_result_1222 = ((_zz_io_result_1213[0] && _zz_io_result_1211[1]) ^ (_zz_io_result_1211[0] && _zz_io_result_1213[1]));
  always @(*) begin
    _zz_io_result_1223[1] = ((_zz_io_result_1213[0] && _zz_io_result_1211[0]) ^ _zz_io_result_1222);
    _zz_io_result_1223[0] = ((_zz_io_result_1213[1] && _zz_io_result_1211[1]) ^ _zz_io_result_1222);
  end

  assign _zz_io_result_1224 = ((_zz_io_result_1214[0] && _zz_io_result_1212[1]) ^ (_zz_io_result_1212[0] && _zz_io_result_1214[1]));
  always @(*) begin
    _zz_io_result_1225[1] = ((_zz_io_result_1214[0] && _zz_io_result_1212[0]) ^ _zz_io_result_1224);
    _zz_io_result_1225[0] = ((_zz_io_result_1214[1] && _zz_io_result_1212[1]) ^ _zz_io_result_1224);
  end

  always @(*) begin
    _zz_io_result_1210[3 : 2] = (_zz_io_result_1223 ^ _zz_io_result_1220);
    _zz_io_result_1210[1 : 0] = (_zz_io_result_1225 ^ _zz_io_result_1220);
  end

  always @(*) begin
    _zz_io_result_1157[7 : 4] = _zz_io_result_1210;
    _zz_io_result_1157[3 : 0] = _zz_io_result_1194;
  end

  assign _zz_io_result_1156 = _zz_io_result_1157;
  always @(*) begin
    _zz_io_result_1227[7] = (_zz_io_result_1156[5] ^ _zz_io_result_1156[3]);
    _zz_io_result_1227[6] = (_zz_io_result_1156[7] ^ _zz_io_result_1156[3]);
    _zz_io_result_1227[5] = (_zz_io_result_1156[6] ^ _zz_io_result_1156[0]);
    _zz_io_result_1227[4] = ((_zz_io_result_1156[7] ^ _zz_io_result_1156[5]) ^ _zz_io_result_1156[3]);
    _zz_io_result_1227[3] = ((((_zz_io_result_1156[7] ^ _zz_io_result_1156[6]) ^ _zz_io_result_1156[5]) ^ _zz_io_result_1156[4]) ^ _zz_io_result_1156[3]);
    _zz_io_result_1227[2] = ((((_zz_io_result_1156[6] ^ _zz_io_result_1156[5]) ^ _zz_io_result_1156[3]) ^ _zz_io_result_1156[2]) ^ _zz_io_result_1156[0]);
    _zz_io_result_1227[1] = ((_zz_io_result_1156[5] ^ _zz_io_result_1156[4]) ^ _zz_io_result_1156[1]);
    _zz_io_result_1227[0] = ((_zz_io_result_1156[6] ^ _zz_io_result_1156[4]) ^ _zz_io_result_1156[1]);
  end

  assign _zz_io_result_1226 = _zz_io_result_1227;
  always @(*) begin
    _zz_io_result_1153[7] = _zz_io_result_1226[7];
    _zz_io_result_1153[6] = (! _zz_io_result_1226[6]);
    _zz_io_result_1153[5] = (! _zz_io_result_1226[5]);
    _zz_io_result_1153[4] = _zz_io_result_1226[4];
    _zz_io_result_1153[3] = _zz_io_result_1226[3];
    _zz_io_result_1153[2] = _zz_io_result_1226[2];
    _zz_io_result_1153[1] = (! _zz_io_result_1226[1]);
    _zz_io_result_1153[0] = (! _zz_io_result_1226[0]);
  end

  assign _zz_io_result_1228 = {_zz_io_result_923,{_zz_io_result_618,{_zz_io_result_313,_zz_io_result_8}}};
  assign _zz_io_result_1233 = {_zz_io_result_1228[127 : 120],{_zz_io_result_1228[87 : 80],{_zz_io_result_1228[47 : 40],{_zz_io_result_1228[7 : 0],{_zz_io_result_1228[95 : 88],{_zz_io_result_1228[55 : 48],{_zz_io_result_1228[15 : 8],{_zz_io_result_1228[103 : 96],{_zz_io_result_1228[63 : 56],{_zz_io_result_1228[23 : 16],{_zz_io_result_1228[111 : 104],{_zz_io_result_1228[71 : 64],{_zz_io_result_1228[31 : 24],{_zz_io_result_1228[119 : 112],{_zz_io_result_1228[79 : 72],_zz_io_result_1228[39 : 32]}}}}}}}}}}}}}}};
  assign _zz_io_result_1229 = _zz_io_result_1233[31 : 0];
  assign _zz_io_result_1230 = _zz_io_result_1233[63 : 32];
  assign _zz_io_result_1231 = _zz_io_result_1233[95 : 64];
  assign _zz_io_result_1232 = _zz_io_result_1233[127 : 96];
  assign _zz_io_result_1235 = {_zz_io_result_1229[7 : 0],_zz_io_result_1229[31 : 8]};
  assign _zz_io_result_1236 = _zz_io_result_1235[23 : 16];
  assign _zz_io_result_1237 = (_zz_io_result_1235[31 : 24] ^ _zz_io_result_1236);
  always @(*) begin
    _zz_io_result_1238[7] = _zz_io_result_1237[6];
    _zz_io_result_1238[6] = _zz_io_result_1237[5];
    _zz_io_result_1238[5] = _zz_io_result_1237[4];
    _zz_io_result_1238[4] = (_zz_io_result_1237[7] ^ _zz_io_result_1237[3]);
    _zz_io_result_1238[3] = (_zz_io_result_1237[7] ^ _zz_io_result_1237[2]);
    _zz_io_result_1238[2] = _zz_io_result_1237[1];
    _zz_io_result_1238[1] = (_zz_io_result_1237[7] ^ _zz_io_result_1237[0]);
    _zz_io_result_1238[0] = _zz_io_result_1237[7];
  end

  always @(*) begin
    _zz_io_result_1234[7 : 0] = ((_zz_io_result_1236 ^ (_zz_io_result_1235[15 : 8] ^ _zz_io_result_1235[7 : 0])) ^ _zz_io_result_1238);
    _zz_io_result_1234[15 : 8] = ((_zz_io_result_1240 ^ (_zz_io_result_1239[15 : 8] ^ _zz_io_result_1239[7 : 0])) ^ _zz_io_result_1242);
    _zz_io_result_1234[23 : 16] = ((_zz_io_result_1244 ^ (_zz_io_result_1243[15 : 8] ^ _zz_io_result_1243[7 : 0])) ^ _zz_io_result_1246);
    _zz_io_result_1234[31 : 24] = ((_zz_io_result_1248 ^ (_zz_io_result_1247[15 : 8] ^ _zz_io_result_1247[7 : 0])) ^ _zz_io_result_1250);
  end

  assign _zz_io_result_1239 = {_zz_io_result_1229[15 : 0],_zz_io_result_1229[31 : 16]};
  assign _zz_io_result_1240 = _zz_io_result_1239[23 : 16];
  assign _zz_io_result_1241 = (_zz_io_result_1239[31 : 24] ^ _zz_io_result_1240);
  always @(*) begin
    _zz_io_result_1242[7] = _zz_io_result_1241[6];
    _zz_io_result_1242[6] = _zz_io_result_1241[5];
    _zz_io_result_1242[5] = _zz_io_result_1241[4];
    _zz_io_result_1242[4] = (_zz_io_result_1241[7] ^ _zz_io_result_1241[3]);
    _zz_io_result_1242[3] = (_zz_io_result_1241[7] ^ _zz_io_result_1241[2]);
    _zz_io_result_1242[2] = _zz_io_result_1241[1];
    _zz_io_result_1242[1] = (_zz_io_result_1241[7] ^ _zz_io_result_1241[0]);
    _zz_io_result_1242[0] = _zz_io_result_1241[7];
  end

  assign _zz_io_result_1243 = {_zz_io_result_1229[23 : 0],_zz_io_result_1229[31 : 24]};
  assign _zz_io_result_1244 = _zz_io_result_1243[23 : 16];
  assign _zz_io_result_1245 = (_zz_io_result_1243[31 : 24] ^ _zz_io_result_1244);
  always @(*) begin
    _zz_io_result_1246[7] = _zz_io_result_1245[6];
    _zz_io_result_1246[6] = _zz_io_result_1245[5];
    _zz_io_result_1246[5] = _zz_io_result_1245[4];
    _zz_io_result_1246[4] = (_zz_io_result_1245[7] ^ _zz_io_result_1245[3]);
    _zz_io_result_1246[3] = (_zz_io_result_1245[7] ^ _zz_io_result_1245[2]);
    _zz_io_result_1246[2] = _zz_io_result_1245[1];
    _zz_io_result_1246[1] = (_zz_io_result_1245[7] ^ _zz_io_result_1245[0]);
    _zz_io_result_1246[0] = _zz_io_result_1245[7];
  end

  assign _zz_io_result_1247 = _zz_io_result_1229[31 : 0];
  assign _zz_io_result_1248 = _zz_io_result_1247[23 : 16];
  assign _zz_io_result_1249 = (_zz_io_result_1247[31 : 24] ^ _zz_io_result_1248);
  always @(*) begin
    _zz_io_result_1250[7] = _zz_io_result_1249[6];
    _zz_io_result_1250[6] = _zz_io_result_1249[5];
    _zz_io_result_1250[5] = _zz_io_result_1249[4];
    _zz_io_result_1250[4] = (_zz_io_result_1249[7] ^ _zz_io_result_1249[3]);
    _zz_io_result_1250[3] = (_zz_io_result_1249[7] ^ _zz_io_result_1249[2]);
    _zz_io_result_1250[2] = _zz_io_result_1249[1];
    _zz_io_result_1250[1] = (_zz_io_result_1249[7] ^ _zz_io_result_1249[0]);
    _zz_io_result_1250[0] = _zz_io_result_1249[7];
  end

  always @(*) begin
    if(io_needMix) begin
      _zz_io_result_4 = _zz_io_result_1234;
    end else begin
      _zz_io_result_4 = _zz_io_result_1229;
    end
  end

  assign _zz_io_result_1252 = {_zz_io_result_1230[7 : 0],_zz_io_result_1230[31 : 8]};
  assign _zz_io_result_1253 = _zz_io_result_1252[23 : 16];
  assign _zz_io_result_1254 = (_zz_io_result_1252[31 : 24] ^ _zz_io_result_1253);
  always @(*) begin
    _zz_io_result_1255[7] = _zz_io_result_1254[6];
    _zz_io_result_1255[6] = _zz_io_result_1254[5];
    _zz_io_result_1255[5] = _zz_io_result_1254[4];
    _zz_io_result_1255[4] = (_zz_io_result_1254[7] ^ _zz_io_result_1254[3]);
    _zz_io_result_1255[3] = (_zz_io_result_1254[7] ^ _zz_io_result_1254[2]);
    _zz_io_result_1255[2] = _zz_io_result_1254[1];
    _zz_io_result_1255[1] = (_zz_io_result_1254[7] ^ _zz_io_result_1254[0]);
    _zz_io_result_1255[0] = _zz_io_result_1254[7];
  end

  always @(*) begin
    _zz_io_result_1251[7 : 0] = ((_zz_io_result_1253 ^ (_zz_io_result_1252[15 : 8] ^ _zz_io_result_1252[7 : 0])) ^ _zz_io_result_1255);
    _zz_io_result_1251[15 : 8] = ((_zz_io_result_1257 ^ (_zz_io_result_1256[15 : 8] ^ _zz_io_result_1256[7 : 0])) ^ _zz_io_result_1259);
    _zz_io_result_1251[23 : 16] = ((_zz_io_result_1261 ^ (_zz_io_result_1260[15 : 8] ^ _zz_io_result_1260[7 : 0])) ^ _zz_io_result_1263);
    _zz_io_result_1251[31 : 24] = ((_zz_io_result_1265 ^ (_zz_io_result_1264[15 : 8] ^ _zz_io_result_1264[7 : 0])) ^ _zz_io_result_1267);
  end

  assign _zz_io_result_1256 = {_zz_io_result_1230[15 : 0],_zz_io_result_1230[31 : 16]};
  assign _zz_io_result_1257 = _zz_io_result_1256[23 : 16];
  assign _zz_io_result_1258 = (_zz_io_result_1256[31 : 24] ^ _zz_io_result_1257);
  always @(*) begin
    _zz_io_result_1259[7] = _zz_io_result_1258[6];
    _zz_io_result_1259[6] = _zz_io_result_1258[5];
    _zz_io_result_1259[5] = _zz_io_result_1258[4];
    _zz_io_result_1259[4] = (_zz_io_result_1258[7] ^ _zz_io_result_1258[3]);
    _zz_io_result_1259[3] = (_zz_io_result_1258[7] ^ _zz_io_result_1258[2]);
    _zz_io_result_1259[2] = _zz_io_result_1258[1];
    _zz_io_result_1259[1] = (_zz_io_result_1258[7] ^ _zz_io_result_1258[0]);
    _zz_io_result_1259[0] = _zz_io_result_1258[7];
  end

  assign _zz_io_result_1260 = {_zz_io_result_1230[23 : 0],_zz_io_result_1230[31 : 24]};
  assign _zz_io_result_1261 = _zz_io_result_1260[23 : 16];
  assign _zz_io_result_1262 = (_zz_io_result_1260[31 : 24] ^ _zz_io_result_1261);
  always @(*) begin
    _zz_io_result_1263[7] = _zz_io_result_1262[6];
    _zz_io_result_1263[6] = _zz_io_result_1262[5];
    _zz_io_result_1263[5] = _zz_io_result_1262[4];
    _zz_io_result_1263[4] = (_zz_io_result_1262[7] ^ _zz_io_result_1262[3]);
    _zz_io_result_1263[3] = (_zz_io_result_1262[7] ^ _zz_io_result_1262[2]);
    _zz_io_result_1263[2] = _zz_io_result_1262[1];
    _zz_io_result_1263[1] = (_zz_io_result_1262[7] ^ _zz_io_result_1262[0]);
    _zz_io_result_1263[0] = _zz_io_result_1262[7];
  end

  assign _zz_io_result_1264 = _zz_io_result_1230[31 : 0];
  assign _zz_io_result_1265 = _zz_io_result_1264[23 : 16];
  assign _zz_io_result_1266 = (_zz_io_result_1264[31 : 24] ^ _zz_io_result_1265);
  always @(*) begin
    _zz_io_result_1267[7] = _zz_io_result_1266[6];
    _zz_io_result_1267[6] = _zz_io_result_1266[5];
    _zz_io_result_1267[5] = _zz_io_result_1266[4];
    _zz_io_result_1267[4] = (_zz_io_result_1266[7] ^ _zz_io_result_1266[3]);
    _zz_io_result_1267[3] = (_zz_io_result_1266[7] ^ _zz_io_result_1266[2]);
    _zz_io_result_1267[2] = _zz_io_result_1266[1];
    _zz_io_result_1267[1] = (_zz_io_result_1266[7] ^ _zz_io_result_1266[0]);
    _zz_io_result_1267[0] = _zz_io_result_1266[7];
  end

  always @(*) begin
    if(io_needMix) begin
      _zz_io_result_5 = _zz_io_result_1251;
    end else begin
      _zz_io_result_5 = _zz_io_result_1230;
    end
  end

  assign _zz_io_result_1269 = {_zz_io_result_1231[7 : 0],_zz_io_result_1231[31 : 8]};
  assign _zz_io_result_1270 = _zz_io_result_1269[23 : 16];
  assign _zz_io_result_1271 = (_zz_io_result_1269[31 : 24] ^ _zz_io_result_1270);
  always @(*) begin
    _zz_io_result_1272[7] = _zz_io_result_1271[6];
    _zz_io_result_1272[6] = _zz_io_result_1271[5];
    _zz_io_result_1272[5] = _zz_io_result_1271[4];
    _zz_io_result_1272[4] = (_zz_io_result_1271[7] ^ _zz_io_result_1271[3]);
    _zz_io_result_1272[3] = (_zz_io_result_1271[7] ^ _zz_io_result_1271[2]);
    _zz_io_result_1272[2] = _zz_io_result_1271[1];
    _zz_io_result_1272[1] = (_zz_io_result_1271[7] ^ _zz_io_result_1271[0]);
    _zz_io_result_1272[0] = _zz_io_result_1271[7];
  end

  always @(*) begin
    _zz_io_result_1268[7 : 0] = ((_zz_io_result_1270 ^ (_zz_io_result_1269[15 : 8] ^ _zz_io_result_1269[7 : 0])) ^ _zz_io_result_1272);
    _zz_io_result_1268[15 : 8] = ((_zz_io_result_1274 ^ (_zz_io_result_1273[15 : 8] ^ _zz_io_result_1273[7 : 0])) ^ _zz_io_result_1276);
    _zz_io_result_1268[23 : 16] = ((_zz_io_result_1278 ^ (_zz_io_result_1277[15 : 8] ^ _zz_io_result_1277[7 : 0])) ^ _zz_io_result_1280);
    _zz_io_result_1268[31 : 24] = ((_zz_io_result_1282 ^ (_zz_io_result_1281[15 : 8] ^ _zz_io_result_1281[7 : 0])) ^ _zz_io_result_1284);
  end

  assign _zz_io_result_1273 = {_zz_io_result_1231[15 : 0],_zz_io_result_1231[31 : 16]};
  assign _zz_io_result_1274 = _zz_io_result_1273[23 : 16];
  assign _zz_io_result_1275 = (_zz_io_result_1273[31 : 24] ^ _zz_io_result_1274);
  always @(*) begin
    _zz_io_result_1276[7] = _zz_io_result_1275[6];
    _zz_io_result_1276[6] = _zz_io_result_1275[5];
    _zz_io_result_1276[5] = _zz_io_result_1275[4];
    _zz_io_result_1276[4] = (_zz_io_result_1275[7] ^ _zz_io_result_1275[3]);
    _zz_io_result_1276[3] = (_zz_io_result_1275[7] ^ _zz_io_result_1275[2]);
    _zz_io_result_1276[2] = _zz_io_result_1275[1];
    _zz_io_result_1276[1] = (_zz_io_result_1275[7] ^ _zz_io_result_1275[0]);
    _zz_io_result_1276[0] = _zz_io_result_1275[7];
  end

  assign _zz_io_result_1277 = {_zz_io_result_1231[23 : 0],_zz_io_result_1231[31 : 24]};
  assign _zz_io_result_1278 = _zz_io_result_1277[23 : 16];
  assign _zz_io_result_1279 = (_zz_io_result_1277[31 : 24] ^ _zz_io_result_1278);
  always @(*) begin
    _zz_io_result_1280[7] = _zz_io_result_1279[6];
    _zz_io_result_1280[6] = _zz_io_result_1279[5];
    _zz_io_result_1280[5] = _zz_io_result_1279[4];
    _zz_io_result_1280[4] = (_zz_io_result_1279[7] ^ _zz_io_result_1279[3]);
    _zz_io_result_1280[3] = (_zz_io_result_1279[7] ^ _zz_io_result_1279[2]);
    _zz_io_result_1280[2] = _zz_io_result_1279[1];
    _zz_io_result_1280[1] = (_zz_io_result_1279[7] ^ _zz_io_result_1279[0]);
    _zz_io_result_1280[0] = _zz_io_result_1279[7];
  end

  assign _zz_io_result_1281 = _zz_io_result_1231[31 : 0];
  assign _zz_io_result_1282 = _zz_io_result_1281[23 : 16];
  assign _zz_io_result_1283 = (_zz_io_result_1281[31 : 24] ^ _zz_io_result_1282);
  always @(*) begin
    _zz_io_result_1284[7] = _zz_io_result_1283[6];
    _zz_io_result_1284[6] = _zz_io_result_1283[5];
    _zz_io_result_1284[5] = _zz_io_result_1283[4];
    _zz_io_result_1284[4] = (_zz_io_result_1283[7] ^ _zz_io_result_1283[3]);
    _zz_io_result_1284[3] = (_zz_io_result_1283[7] ^ _zz_io_result_1283[2]);
    _zz_io_result_1284[2] = _zz_io_result_1283[1];
    _zz_io_result_1284[1] = (_zz_io_result_1283[7] ^ _zz_io_result_1283[0]);
    _zz_io_result_1284[0] = _zz_io_result_1283[7];
  end

  always @(*) begin
    if(io_needMix) begin
      _zz_io_result_6 = _zz_io_result_1268;
    end else begin
      _zz_io_result_6 = _zz_io_result_1231;
    end
  end

  assign _zz_io_result_1286 = {_zz_io_result_1232[7 : 0],_zz_io_result_1232[31 : 8]};
  assign _zz_io_result_1287 = _zz_io_result_1286[23 : 16];
  assign _zz_io_result_1288 = (_zz_io_result_1286[31 : 24] ^ _zz_io_result_1287);
  always @(*) begin
    _zz_io_result_1289[7] = _zz_io_result_1288[6];
    _zz_io_result_1289[6] = _zz_io_result_1288[5];
    _zz_io_result_1289[5] = _zz_io_result_1288[4];
    _zz_io_result_1289[4] = (_zz_io_result_1288[7] ^ _zz_io_result_1288[3]);
    _zz_io_result_1289[3] = (_zz_io_result_1288[7] ^ _zz_io_result_1288[2]);
    _zz_io_result_1289[2] = _zz_io_result_1288[1];
    _zz_io_result_1289[1] = (_zz_io_result_1288[7] ^ _zz_io_result_1288[0]);
    _zz_io_result_1289[0] = _zz_io_result_1288[7];
  end

  always @(*) begin
    _zz_io_result_1285[7 : 0] = ((_zz_io_result_1287 ^ (_zz_io_result_1286[15 : 8] ^ _zz_io_result_1286[7 : 0])) ^ _zz_io_result_1289);
    _zz_io_result_1285[15 : 8] = ((_zz_io_result_1291 ^ (_zz_io_result_1290[15 : 8] ^ _zz_io_result_1290[7 : 0])) ^ _zz_io_result_1293);
    _zz_io_result_1285[23 : 16] = ((_zz_io_result_1295 ^ (_zz_io_result_1294[15 : 8] ^ _zz_io_result_1294[7 : 0])) ^ _zz_io_result_1297);
    _zz_io_result_1285[31 : 24] = ((_zz_io_result_1299 ^ (_zz_io_result_1298[15 : 8] ^ _zz_io_result_1298[7 : 0])) ^ _zz_io_result_1301);
  end

  assign _zz_io_result_1290 = {_zz_io_result_1232[15 : 0],_zz_io_result_1232[31 : 16]};
  assign _zz_io_result_1291 = _zz_io_result_1290[23 : 16];
  assign _zz_io_result_1292 = (_zz_io_result_1290[31 : 24] ^ _zz_io_result_1291);
  always @(*) begin
    _zz_io_result_1293[7] = _zz_io_result_1292[6];
    _zz_io_result_1293[6] = _zz_io_result_1292[5];
    _zz_io_result_1293[5] = _zz_io_result_1292[4];
    _zz_io_result_1293[4] = (_zz_io_result_1292[7] ^ _zz_io_result_1292[3]);
    _zz_io_result_1293[3] = (_zz_io_result_1292[7] ^ _zz_io_result_1292[2]);
    _zz_io_result_1293[2] = _zz_io_result_1292[1];
    _zz_io_result_1293[1] = (_zz_io_result_1292[7] ^ _zz_io_result_1292[0]);
    _zz_io_result_1293[0] = _zz_io_result_1292[7];
  end

  assign _zz_io_result_1294 = {_zz_io_result_1232[23 : 0],_zz_io_result_1232[31 : 24]};
  assign _zz_io_result_1295 = _zz_io_result_1294[23 : 16];
  assign _zz_io_result_1296 = (_zz_io_result_1294[31 : 24] ^ _zz_io_result_1295);
  always @(*) begin
    _zz_io_result_1297[7] = _zz_io_result_1296[6];
    _zz_io_result_1297[6] = _zz_io_result_1296[5];
    _zz_io_result_1297[5] = _zz_io_result_1296[4];
    _zz_io_result_1297[4] = (_zz_io_result_1296[7] ^ _zz_io_result_1296[3]);
    _zz_io_result_1297[3] = (_zz_io_result_1296[7] ^ _zz_io_result_1296[2]);
    _zz_io_result_1297[2] = _zz_io_result_1296[1];
    _zz_io_result_1297[1] = (_zz_io_result_1296[7] ^ _zz_io_result_1296[0]);
    _zz_io_result_1297[0] = _zz_io_result_1296[7];
  end

  assign _zz_io_result_1298 = _zz_io_result_1232[31 : 0];
  assign _zz_io_result_1299 = _zz_io_result_1298[23 : 16];
  assign _zz_io_result_1300 = (_zz_io_result_1298[31 : 24] ^ _zz_io_result_1299);
  always @(*) begin
    _zz_io_result_1301[7] = _zz_io_result_1300[6];
    _zz_io_result_1301[6] = _zz_io_result_1300[5];
    _zz_io_result_1301[5] = _zz_io_result_1300[4];
    _zz_io_result_1301[4] = (_zz_io_result_1300[7] ^ _zz_io_result_1300[3]);
    _zz_io_result_1301[3] = (_zz_io_result_1300[7] ^ _zz_io_result_1300[2]);
    _zz_io_result_1301[2] = _zz_io_result_1300[1];
    _zz_io_result_1301[1] = (_zz_io_result_1300[7] ^ _zz_io_result_1300[0]);
    _zz_io_result_1301[0] = _zz_io_result_1300[7];
  end

  always @(*) begin
    if(io_needMix) begin
      _zz_io_result_7 = _zz_io_result_1285;
    end else begin
      _zz_io_result_7 = _zz_io_result_1232;
    end
  end

  assign io_result = {_zz_io_result_7,{_zz_io_result_6,{_zz_io_result_5,_zz_io_result_4}}};

endmodule
